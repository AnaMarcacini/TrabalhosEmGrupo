<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-92.2026,38.2799,300.387,-164.198</PageViewport>
<gate>
<ID>965</ID>
<type>DA_FROM</type>
<position>85.5,-39.5</position>
<input>
<ID>IN_0</ID>738 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D3_IR</lparam></gate>
<gate>
<ID>193</ID>
<type>AA_MUX_2x1</type>
<position>94,-85</position>
<input>
<ID>IN_0</ID>760 </input>
<input>
<ID>IN_1</ID>761 </input>
<output>
<ID>OUT</ID>759 </output>
<input>
<ID>SEL_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>966</ID>
<type>DA_FROM</type>
<position>88.5,-70</position>
<input>
<ID>IN_0</ID>758 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D7_IR</lparam></gate>
<gate>
<ID>194</ID>
<type>AA_MUX_2x1</type>
<position>94.5,-90</position>
<input>
<ID>IN_0</ID>770 </input>
<input>
<ID>IN_1</ID>762 </input>
<output>
<ID>OUT</ID>769 </output>
<input>
<ID>SEL_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1</ID>
<type>DE_TO</type>
<position>32,-6</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA0</lparam></gate>
<gate>
<ID>967</ID>
<type>DA_FROM</type>
<position>76.5,-53</position>
<input>
<ID>IN_0</ID>749 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D4_IR</lparam></gate>
<gate>
<ID>195</ID>
<type>AA_MUX_2x1</type>
<position>94.5,-95.5</position>
<input>
<ID>IN_0</ID>768 </input>
<input>
<ID>IN_1</ID>763 </input>
<output>
<ID>OUT</ID>767 </output>
<input>
<ID>SEL_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2</ID>
<type>DE_TO</type>
<position>32,-19</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA1</lparam></gate>
<gate>
<ID>968</ID>
<type>DA_FROM</type>
<position>86,-59</position>
<input>
<ID>IN_0</ID>752 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D5_IR</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_MUX_2x1</type>
<position>95,-101.5</position>
<input>
<ID>IN_0</ID>765 </input>
<input>
<ID>IN_1</ID>764 </input>
<output>
<ID>OUT</ID>766 </output>
<input>
<ID>SEL_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>DE_TO</type>
<position>32,-32</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA2</lparam></gate>
<gate>
<ID>4</ID>
<type>DE_TO</type>
<position>32,-45</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA3</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_AND4</type>
<position>81,3</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>80 </input>
<input>
<ID>IN_2</ID>81 </input>
<input>
<ID>IN_3</ID>86 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>5</ID>
<type>DE_TO</type>
<position>32,-58</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA4</lparam></gate>
<gate>
<ID>971</ID>
<type>DA_FROM</type>
<position>88,-63.5</position>
<input>
<ID>IN_0</ID>754 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D6_IR</lparam></gate>
<gate>
<ID>6</ID>
<type>DE_TO</type>
<position>32,-70</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA5</lparam></gate>
<gate>
<ID>972</ID>
<type>DA_FROM</type>
<position>87,-100</position>
<input>
<ID>IN_0</ID>764 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D11_IR</lparam></gate>
<gate>
<ID>7</ID>
<type>DE_TO</type>
<position>32,-83</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA6</lparam></gate>
<gate>
<ID>973</ID>
<type>DA_FROM</type>
<position>81.5,-83</position>
<input>
<ID>IN_0</ID>761 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D8_IR</lparam></gate>
<gate>
<ID>8</ID>
<type>DE_TO</type>
<position>32,-96</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA7</lparam></gate>
<gate>
<ID>974</ID>
<type>DA_FROM</type>
<position>86.5,-87.5</position>
<input>
<ID>IN_0</ID>762 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D9_IR</lparam></gate>
<gate>
<ID>202</ID>
<type>DA_FROM</type>
<position>72.5,6</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_IR</lparam></gate>
<gate>
<ID>9</ID>
<type>DE_TO</type>
<position>32,-109</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA8</lparam></gate>
<gate>
<ID>975</ID>
<type>DA_FROM</type>
<position>89,-93.5</position>
<input>
<ID>IN_0</ID>763 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D10_IR</lparam></gate>
<gate>
<ID>203</ID>
<type>DA_FROM</type>
<position>64.5,3.5</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D14_IR</lparam></gate>
<gate>
<ID>10</ID>
<type>DE_TO</type>
<position>32,-122</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA9</lparam></gate>
<gate>
<ID>11</ID>
<type>DE_TO</type>
<position>32,-135</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA10</lparam></gate>
<gate>
<ID>12</ID>
<type>DE_TO</type>
<position>32,-148</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA11</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>30.5,31</position>
<gparam>LABEL_TEXT PROCESSADOR BIP IMT - MAUA 2022</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>44</ID>
<type>AE_DFF_LOW_NT</type>
<position>22,-6</position>
<input>
<ID>IN_0</ID>43 </input>
<output>
<ID>OUT_0</ID>13 </output>
<input>
<ID>clear</ID>74 </input>
<input>
<ID>clock</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_DFF_LOW_NT</type>
<position>22,-19</position>
<input>
<ID>IN_0</ID>44 </input>
<output>
<ID>OUT_0</ID>14 </output>
<input>
<ID>clear</ID>74 </input>
<input>
<ID>clock</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>46</ID>
<type>AE_DFF_LOW_NT</type>
<position>22,-32</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>15 </output>
<input>
<ID>clear</ID>74 </input>
<input>
<ID>clock</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>47</ID>
<type>AE_DFF_LOW_NT</type>
<position>22,-45</position>
<input>
<ID>IN_0</ID>46 </input>
<output>
<ID>OUT_0</ID>16 </output>
<input>
<ID>clear</ID>74 </input>
<input>
<ID>clock</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>48</ID>
<type>AE_DFF_LOW_NT</type>
<position>22,-58</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>19 </output>
<input>
<ID>clear</ID>74 </input>
<input>
<ID>clock</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>49</ID>
<type>AE_DFF_LOW_NT</type>
<position>22,-70</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>20 </output>
<input>
<ID>clear</ID>74 </input>
<input>
<ID>clock</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>50</ID>
<type>AE_DFF_LOW_NT</type>
<position>22,-83</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>21 </output>
<input>
<ID>clear</ID>74 </input>
<input>
<ID>clock</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>51</ID>
<type>AE_DFF_LOW_NT</type>
<position>22,-96</position>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT_0</ID>22 </output>
<input>
<ID>clear</ID>74 </input>
<input>
<ID>clock</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>52</ID>
<type>AE_DFF_LOW_NT</type>
<position>22,-109</position>
<input>
<ID>IN_0</ID>51 </input>
<output>
<ID>OUT_0</ID>26 </output>
<input>
<ID>clear</ID>74 </input>
<input>
<ID>clock</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>53</ID>
<type>AE_DFF_LOW_NT</type>
<position>22,-122</position>
<input>
<ID>IN_0</ID>52 </input>
<output>
<ID>OUT_0</ID>27 </output>
<input>
<ID>clear</ID>74 </input>
<input>
<ID>clock</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>54</ID>
<type>AE_DFF_LOW_NT</type>
<position>22,-135</position>
<input>
<ID>IN_0</ID>53 </input>
<output>
<ID>OUT_0</ID>28 </output>
<input>
<ID>clear</ID>74 </input>
<input>
<ID>clock</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>55</ID>
<type>AE_DFF_LOW_NT</type>
<position>22,-148</position>
<input>
<ID>IN_0</ID>54 </input>
<output>
<ID>OUT_0</ID>29 </output>
<input>
<ID>clear</ID>74 </input>
<input>
<ID>clock</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>57</ID>
<type>AE_FULLADDER_4BIT</type>
<position>61,-31</position>
<input>
<ID>IN_0</ID>825 </input>
<input>
<ID>IN_1</ID>25 </input>
<input>
<ID>IN_2</ID>25 </input>
<input>
<ID>IN_3</ID>25 </input>
<input>
<ID>IN_B_0</ID>13 </input>
<input>
<ID>IN_B_1</ID>14 </input>
<input>
<ID>IN_B_2</ID>15 </input>
<input>
<ID>IN_B_3</ID>16 </input>
<output>
<ID>OUT_0</ID>118 </output>
<output>
<ID>OUT_1</ID>125 </output>
<output>
<ID>OUT_2</ID>734 </output>
<output>
<ID>OUT_3</ID>737 </output>
<input>
<ID>carry_in</ID>12 </input>
<output>
<ID>carry_out</ID>10 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>60</ID>
<type>AE_FULLADDER_4BIT</type>
<position>61,-62</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>23 </input>
<input>
<ID>IN_2</ID>23 </input>
<input>
<ID>IN_3</ID>23 </input>
<input>
<ID>IN_B_0</ID>19 </input>
<input>
<ID>IN_B_1</ID>20 </input>
<input>
<ID>IN_B_2</ID>21 </input>
<input>
<ID>IN_B_3</ID>22 </input>
<output>
<ID>OUT_0</ID>744 </output>
<output>
<ID>OUT_1</ID>751 </output>
<output>
<ID>OUT_2</ID>755 </output>
<output>
<ID>OUT_3</ID>757 </output>
<input>
<ID>carry_in</ID>10 </input>
<output>
<ID>carry_out</ID>11 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>61</ID>
<type>AE_FULLADDER_4BIT</type>
<position>61,-91</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>30 </input>
<input>
<ID>IN_2</ID>30 </input>
<input>
<ID>IN_3</ID>30 </input>
<input>
<ID>IN_B_0</ID>26 </input>
<input>
<ID>IN_B_1</ID>27 </input>
<input>
<ID>IN_B_2</ID>28 </input>
<input>
<ID>IN_B_3</ID>29 </input>
<output>
<ID>OUT_0</ID>760 </output>
<output>
<ID>OUT_1</ID>770 </output>
<output>
<ID>OUT_2</ID>768 </output>
<output>
<ID>OUT_3</ID>765 </output>
<input>
<ID>carry_in</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>63</ID>
<type>FF_GND</type>
<position>62.5,-20</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>67</ID>
<type>FF_GND</type>
<position>56,-39</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>69</ID>
<type>FF_GND</type>
<position>56,-68.5</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>71</ID>
<type>FF_GND</type>
<position>56,-99</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>75</ID>
<type>DE_TO</type>
<position>102.5,-30.5</position>
<input>
<ID>IN_0</ID>123 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA1</lparam></gate>
<gate>
<ID>76</ID>
<type>DE_TO</type>
<position>102,-36</position>
<input>
<ID>IN_0</ID>733 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA2</lparam></gate>
<gate>
<ID>77</ID>
<type>DE_TO</type>
<position>102,-40.5</position>
<input>
<ID>IN_0</ID>736 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA3</lparam></gate>
<gate>
<ID>849</ID>
<type>AA_LABEL</type>
<position>95,-114</position>
<gparam>LABEL_TEXT Sinais de Controle</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>DE_TO</type>
<position>104,-55.5</position>
<input>
<ID>IN_0</ID>743 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA4</lparam></gate>
<gate>
<ID>79</ID>
<type>DE_TO</type>
<position>103.5,-60.5</position>
<input>
<ID>IN_0</ID>750 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA5</lparam></gate>
<gate>
<ID>851</ID>
<type>AA_LABEL</type>
<position>75.5,-121.5</position>
<gparam>LABEL_TEXT RESET</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>DE_TO</type>
<position>103.5,-65.5</position>
<input>
<ID>IN_0</ID>753 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA6</lparam></gate>
<gate>
<ID>852</ID>
<type>AA_LABEL</type>
<position>75.5,-126.5</position>
<gparam>LABEL_TEXT WR_PC</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>DE_TO</type>
<position>104,-71.5</position>
<input>
<ID>IN_0</ID>756 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA7</lparam></gate>
<gate>
<ID>853</ID>
<type>AA_LABEL</type>
<position>76,-132</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>DE_TO</type>
<position>101,-84.5</position>
<input>
<ID>IN_0</ID>759 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA8</lparam></gate>
<gate>
<ID>83</ID>
<type>DE_TO</type>
<position>101,-90</position>
<input>
<ID>IN_0</ID>769 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA9</lparam></gate>
<gate>
<ID>84</ID>
<type>DE_TO</type>
<position>102.5,-96</position>
<input>
<ID>IN_0</ID>767 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA10</lparam></gate>
<gate>
<ID>85</ID>
<type>DE_TO</type>
<position>103,-101.5</position>
<input>
<ID>IN_0</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA11</lparam></gate>
<gate>
<ID>87</ID>
<type>DA_FROM</type>
<position>13,-4</position>
<input>
<ID>IN_0</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA0</lparam></gate>
<gate>
<ID>88</ID>
<type>DA_FROM</type>
<position>13,-17</position>
<input>
<ID>IN_0</ID>44 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA1</lparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>13,-30</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA2</lparam></gate>
<gate>
<ID>90</ID>
<type>DA_FROM</type>
<position>13,-43</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA3</lparam></gate>
<gate>
<ID>93</ID>
<type>DA_FROM</type>
<position>13,-56</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA4</lparam></gate>
<gate>
<ID>94</ID>
<type>DA_FROM</type>
<position>13,-68</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA5</lparam></gate>
<gate>
<ID>95</ID>
<type>DA_FROM</type>
<position>13,-81</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA6</lparam></gate>
<gate>
<ID>96</ID>
<type>DA_FROM</type>
<position>13,-94</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA7</lparam></gate>
<gate>
<ID>97</ID>
<type>DA_FROM</type>
<position>13,-107</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA8</lparam></gate>
<gate>
<ID>98</ID>
<type>DA_FROM</type>
<position>13,-120</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA9</lparam></gate>
<gate>
<ID>99</ID>
<type>DA_FROM</type>
<position>13,-133</position>
<input>
<ID>IN_0</ID>53 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA10</lparam></gate>
<gate>
<ID>100</ID>
<type>DA_FROM</type>
<position>13,-146</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA11</lparam></gate>
<gate>
<ID>102</ID>
<type>DA_FROM</type>
<position>-8,-6.5</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>24,8</position>
<gparam>LABEL_TEXT Contador de Programa - PC</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>27.5,19</position>
<gparam>LABEL_TEXT Prof.  Angelo Zanini / Nuncio Perrella</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>124</ID>
<type>DA_FROM</type>
<position>53.5,-33</position>
<input>
<ID>IN_0</ID>825 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WR_PC</lparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>-8,-11.5</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RESET</lparam></gate>
<gate>
<ID>136</ID>
<type>DA_FROM</type>
<position>84,-15</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D0_IR</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_MUX_2x1</type>
<position>94,-24.5</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>89 </output>
<input>
<ID>SEL_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>AA_MUX_2x1</type>
<position>94.5,-29.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>123 </output>
<input>
<ID>SEL_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_MUX_2x1</type>
<position>94.5,-35</position>
<input>
<ID>IN_0</ID>734 </input>
<input>
<ID>IN_1</ID>735 </input>
<output>
<ID>OUT</ID>733 </output>
<input>
<ID>SEL_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>927</ID>
<type>DA_FROM</type>
<position>64.5,0.5</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D13_IR</lparam></gate>
<gate>
<ID>928</ID>
<type>DA_FROM</type>
<position>64.5,-2.5</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D12_IR</lparam></gate>
<gate>
<ID>932</ID>
<type>AE_SMALL_INVERTER</type>
<position>73,3.5</position>
<input>
<ID>IN_0</ID>79 </input>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>933</ID>
<type>AE_SMALL_INVERTER</type>
<position>73,1</position>
<input>
<ID>IN_0</ID>82 </input>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>934</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-2.5</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>936</ID>
<type>DE_TO</type>
<position>94,3</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Saida</lparam></gate>
<gate>
<ID>939</ID>
<type>DE_TO</type>
<position>102,-24.5</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PA0</lparam></gate>
<gate>
<ID>944</ID>
<type>AA_MUX_2x1</type>
<position>139.5,-59.5</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>122 </output>
<input>
<ID>SEL_0</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>947</ID>
<type>AA_TOGGLE</type>
<position>137.5,-49</position>
<output>
<ID>OUT_0</ID>119 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>952</ID>
<type>FF_GND</type>
<position>131,-62.5</position>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>959</ID>
<type>EE_VDD</type>
<position>131.5,-55</position>
<output>
<ID>OUT_0</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_MUX_2x1</type>
<position>95,-41</position>
<input>
<ID>IN_0</ID>737 </input>
<input>
<ID>IN_1</ID>738 </input>
<output>
<ID>OUT</ID>736 </output>
<input>
<ID>SEL_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_MUX_2x1</type>
<position>94.5,-55.5</position>
<input>
<ID>IN_0</ID>744 </input>
<input>
<ID>IN_1</ID>749 </input>
<output>
<ID>OUT</ID>743 </output>
<input>
<ID>SEL_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>962</ID>
<type>GA_LED</type>
<position>149,-60</position>
<input>
<ID>N_in0</ID>122 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>AA_MUX_2x1</type>
<position>95,-60.5</position>
<input>
<ID>IN_0</ID>751 </input>
<input>
<ID>IN_1</ID>752 </input>
<output>
<ID>OUT</ID>750 </output>
<input>
<ID>SEL_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>963</ID>
<type>DA_FROM</type>
<position>85,-28</position>
<input>
<ID>IN_0</ID>126 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D1_IR</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_MUX_2x1</type>
<position>95,-66</position>
<input>
<ID>IN_0</ID>755 </input>
<input>
<ID>IN_1</ID>754 </input>
<output>
<ID>OUT</ID>753 </output>
<input>
<ID>SEL_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>964</ID>
<type>DA_FROM</type>
<position>87,-33</position>
<input>
<ID>IN_0</ID>735 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID D2_IR</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_MUX_2x1</type>
<position>95.5,-72</position>
<input>
<ID>IN_0</ID>757 </input>
<input>
<ID>IN_1</ID>758 </input>
<output>
<ID>OUT</ID>756 </output>
<input>
<ID>SEL_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-54,60,-39</points>
<connection>
<GID>60</GID>
<name>carry_in</name></connection>
<connection>
<GID>57</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-83,60,-70</points>
<connection>
<GID>60</GID>
<name>carry_out</name></connection>
<connection>
<GID>61</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>60,-23,60,-19</points>
<connection>
<GID>57</GID>
<name>carry_in</name></connection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>60,-19,62.5,-19</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<intersection>60 1</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-26,41,-4</points>
<intersection>-26 1</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-26,57,-26</points>
<connection>
<GID>57</GID>
<name>IN_B_0</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-4,41,-4</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>28 3</intersection>
<intersection>41 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-6,28,-4</points>
<intersection>-6 4</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28,-6,30,-6</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>28 3</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-27,40,-17</points>
<intersection>-27 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-27,57,-27</points>
<connection>
<GID>57</GID>
<name>IN_B_1</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-17,40,-17</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>28 3</intersection>
<intersection>40 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-19,28,-17</points>
<intersection>-19 4</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28,-19,30,-19</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>28 3</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-30,39,-28</points>
<intersection>-30 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-28,57,-28</points>
<connection>
<GID>57</GID>
<name>IN_B_2</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-30,39,-30</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>28 3</intersection>
<intersection>39 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-32,28,-30</points>
<intersection>-32 4</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28,-32,30,-32</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>28 3</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-43,41,-29</points>
<intersection>-43 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-29,57,-29</points>
<connection>
<GID>57</GID>
<name>IN_B_3</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-43,41,-43</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>28 3</intersection>
<intersection>41 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-45,28,-43</points>
<intersection>-45 4</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28,-45,30,-45</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>28 3</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-57,41,-56</points>
<intersection>-57 1</intersection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-57,57,-57</points>
<connection>
<GID>60</GID>
<name>IN_B_0</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-56,41,-56</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>28 3</intersection>
<intersection>41 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-58,28,-56</points>
<intersection>-58 4</intersection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28,-58,30,-58</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>28 3</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-68,41,-58</points>
<intersection>-68 2</intersection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-58,57,-58</points>
<connection>
<GID>60</GID>
<name>IN_B_1</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-68,41,-68</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>28 3</intersection>
<intersection>41 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-70,28,-68</points>
<intersection>-70 4</intersection>
<intersection>-68 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28,-70,30,-70</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>28 3</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-81,44,-59</points>
<intersection>-81 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-59,57,-59</points>
<connection>
<GID>60</GID>
<name>IN_B_2</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-81,44,-81</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>28 3</intersection>
<intersection>44 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-83,28,-81</points>
<intersection>-83 4</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28,-83,30,-83</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>28 3</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-94,47,-60</points>
<intersection>-94 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-60,57,-60</points>
<connection>
<GID>60</GID>
<name>IN_B_3</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-94,47,-94</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>28 3</intersection>
<intersection>47 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-96,28,-94</points>
<intersection>-96 4</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28,-96,30,-96</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>28 3</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-67.5,56,-64</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>-67 1</intersection>
<intersection>-66 7</intersection>
<intersection>-65 6</intersection>
<intersection>-64 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-67,57,-67</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>56,-64,57,-64</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>56,-65,57,-65</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>56,-66,57,-66</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-38,56,-34</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>-36 4</intersection>
<intersection>-35 6</intersection>
<intersection>-34 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>56,-36,57,-36</points>
<connection>
<GID>57</GID>
<name>IN_3</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>56,-34,57,-34</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>56,-35,57,-35</points>
<connection>
<GID>57</GID>
<name>IN_2</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-107,48,-86</points>
<intersection>-107 2</intersection>
<intersection>-86 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-86,57,-86</points>
<connection>
<GID>61</GID>
<name>IN_B_0</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-107,48,-107</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>28 3</intersection>
<intersection>48 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-109,28,-107</points>
<intersection>-109 4</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28,-109,30,-109</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>28 3</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-120,49,-87</points>
<intersection>-120 2</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-87,57,-87</points>
<connection>
<GID>61</GID>
<name>IN_B_1</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-120,49,-120</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>28 3</intersection>
<intersection>49 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-122,28,-120</points>
<intersection>-122 4</intersection>
<intersection>-120 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28,-122,30,-122</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>28 3</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-133,50,-88</points>
<intersection>-133 2</intersection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-88,57,-88</points>
<connection>
<GID>61</GID>
<name>IN_B_2</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-133,50,-133</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>28 3</intersection>
<intersection>50 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-135,28,-133</points>
<intersection>-135 4</intersection>
<intersection>-133 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28,-135,30,-135</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>28 3</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-146,51,-89</points>
<intersection>-146 2</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-89,57,-89</points>
<connection>
<GID>61</GID>
<name>IN_B_3</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-146,51,-146</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>28 3</intersection>
<intersection>51 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-148,28,-146</points>
<intersection>-148 4</intersection>
<intersection>-146 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28,-148,30,-148</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>28 3</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-98,56,-93</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>-96 1</intersection>
<intersection>-95 5</intersection>
<intersection>-94 4</intersection>
<intersection>-93 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-96,57,-96</points>
<connection>
<GID>61</GID>
<name>IN_3</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>56,-94,57,-94</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>56,-95,57,-95</points>
<connection>
<GID>61</GID>
<name>IN_2</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>56,-93,57,-93</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-4,19,-4</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-17,19,-17</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<connection>
<GID>88</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-30,19,-30</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<connection>
<GID>89</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-43,19,-43</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<connection>
<GID>90</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-56,19,-56</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<connection>
<GID>93</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-68,19,-68</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-81,19,-81</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<connection>
<GID>95</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-94,19,-94</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<connection>
<GID>96</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-107,19,-107</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<connection>
<GID>97</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-120,19,-120</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<connection>
<GID>98</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>825</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,-33,57,-33</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<connection>
<GID>124</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-133,19,-133</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<connection>
<GID>99</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-146,19,-146</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<connection>
<GID>100</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,-6.5,19,-6.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>0 3</intersection>
<intersection>19 26</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>0,-149,0,-6.5</points>
<intersection>-149 25</intersection>
<intersection>-136 23</intersection>
<intersection>-123 21</intersection>
<intersection>-110 19</intersection>
<intersection>-97 17</intersection>
<intersection>-84 15</intersection>
<intersection>-71 13</intersection>
<intersection>-59 11</intersection>
<intersection>-46 9</intersection>
<intersection>-33 7</intersection>
<intersection>-20 4</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>0,-20,19,-20</points>
<connection>
<GID>45</GID>
<name>clock</name></connection>
<intersection>0 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>0,-33,19,-33</points>
<connection>
<GID>46</GID>
<name>clock</name></connection>
<intersection>0 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>0,-46,19,-46</points>
<connection>
<GID>47</GID>
<name>clock</name></connection>
<intersection>0 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>0,-59,19,-59</points>
<connection>
<GID>48</GID>
<name>clock</name></connection>
<intersection>0 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>0,-71,19,-71</points>
<connection>
<GID>49</GID>
<name>clock</name></connection>
<intersection>0 3</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>0,-84,19,-84</points>
<connection>
<GID>50</GID>
<name>clock</name></connection>
<intersection>0 3</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>0,-97,19,-97</points>
<connection>
<GID>51</GID>
<name>clock</name></connection>
<intersection>0 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>0,-110,19,-110</points>
<connection>
<GID>52</GID>
<name>clock</name></connection>
<intersection>0 3</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>0,-123,19,-123</points>
<connection>
<GID>53</GID>
<name>clock</name></connection>
<intersection>0 3</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>0,-136,19,-136</points>
<connection>
<GID>54</GID>
<name>clock</name></connection>
<intersection>0 3</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>0,-149,19,-149</points>
<connection>
<GID>55</GID>
<name>clock</name></connection>
<intersection>0 3</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>19,-7,19,-6.5</points>
<connection>
<GID>44</GID>
<name>clock</name></connection>
<intersection>-6.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,-11.5,22,-11.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-3 2</intersection>
<intersection>22 41</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-3,-153,-3,-11.5</points>
<intersection>-153 29</intersection>
<intersection>-140 28</intersection>
<intersection>-127 26</intersection>
<intersection>-114 24</intersection>
<intersection>-101 22</intersection>
<intersection>-88 20</intersection>
<intersection>-75 18</intersection>
<intersection>-63 16</intersection>
<intersection>-50 14</intersection>
<intersection>-37 12</intersection>
<intersection>-24 10</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-3,-24,22,-24</points>
<intersection>-3 2</intersection>
<intersection>22 40</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-3,-37,22,-37</points>
<intersection>-3 2</intersection>
<intersection>22 39</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-3,-50,22,-50</points>
<intersection>-3 2</intersection>
<intersection>22 38</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-3,-63,22,-63</points>
<intersection>-3 2</intersection>
<intersection>22 37</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-3,-75,22,-75</points>
<intersection>-3 2</intersection>
<intersection>22 36</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-3,-88,22,-88</points>
<intersection>-3 2</intersection>
<intersection>22 35</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-3,-101,22,-101</points>
<intersection>-3 2</intersection>
<intersection>22 34</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>-3,-114,22,-114</points>
<intersection>-3 2</intersection>
<intersection>22 33</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-3,-127,22,-127</points>
<intersection>-3 2</intersection>
<intersection>22 32</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-3,-140,22,-140</points>
<intersection>-3 2</intersection>
<intersection>22 31</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>-3,-153,22,-153</points>
<intersection>-3 2</intersection>
<intersection>22 30</intersection></hsegment>
<vsegment>
<ID>30</ID>
<points>22,-153,22,-152</points>
<connection>
<GID>55</GID>
<name>clear</name></connection>
<intersection>-153 29</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>22,-140,22,-139</points>
<connection>
<GID>54</GID>
<name>clear</name></connection>
<intersection>-140 28</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>22,-127,22,-126</points>
<connection>
<GID>53</GID>
<name>clear</name></connection>
<intersection>-127 26</intersection></vsegment>
<vsegment>
<ID>33</ID>
<points>22,-114,22,-113</points>
<connection>
<GID>52</GID>
<name>clear</name></connection>
<intersection>-114 24</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>22,-101,22,-100</points>
<connection>
<GID>51</GID>
<name>clear</name></connection>
<intersection>-101 22</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>22,-88,22,-87</points>
<connection>
<GID>50</GID>
<name>clear</name></connection>
<intersection>-88 20</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>22,-75,22,-74</points>
<connection>
<GID>49</GID>
<name>clear</name></connection>
<intersection>-75 18</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>22,-63,22,-62</points>
<connection>
<GID>48</GID>
<name>clear</name></connection>
<intersection>-63 16</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>22,-50,22,-49</points>
<connection>
<GID>47</GID>
<name>clear</name></connection>
<intersection>-50 14</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>22,-37,22,-36</points>
<connection>
<GID>46</GID>
<name>clear</name></connection>
<intersection>-37 12</intersection></vsegment>
<vsegment>
<ID>40</ID>
<points>22,-24,22,-23</points>
<connection>
<GID>45</GID>
<name>clear</name></connection>
<intersection>-24 10</intersection></vsegment>
<vsegment>
<ID>41</ID>
<points>22,-11.5,22,-10</points>
<connection>
<GID>44</GID>
<name>clear</name></connection>
<intersection>-11.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,6,78,6</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<connection>
<GID>202</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>66.5,3.5,71,3.5</points>
<connection>
<GID>932</GID>
<name>IN_0</name></connection>
<connection>
<GID>203</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,3.5,76.5,4</points>
<intersection>3.5 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,4,78,4</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,3.5,76.5,3.5</points>
<connection>
<GID>932</GID>
<name>OUT_0</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,1,76.5,2</points>
<intersection>1 2</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,2,78,2</points>
<connection>
<GID>198</GID>
<name>IN_2</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,1,76.5,1</points>
<connection>
<GID>933</GID>
<name>OUT_0</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,0.5,68.5,1</points>
<intersection>0.5 2</intersection>
<intersection>1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,1,71,1</points>
<connection>
<GID>933</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66.5,0.5,68.5,0.5</points>
<connection>
<GID>927</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>66.5,-2.5,70.5,-2.5</points>
<connection>
<GID>928</GID>
<name>IN_0</name></connection>
<intersection>70.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>70.5,-2.5,70.5,-2.5</points>
<connection>
<GID>934</GID>
<name>IN_0</name></connection>
<intersection>-2.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-2.5,76,0</points>
<intersection>-2.5 2</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,0,78,0</points>
<connection>
<GID>198</GID>
<name>IN_3</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-2.5,76,-2.5</points>
<connection>
<GID>934</GID>
<name>OUT_0</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,3,94,3</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<connection>
<GID>936</GID>
<name>IN_0</name></connection>
<intersection>94 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>94,-82.5,94,3</points>
<connection>
<GID>144</GID>
<name>SEL_0</name></connection>
<intersection>-82.5 12</intersection>
<intersection>-69.5 11</intersection>
<intersection>-63.5 26</intersection>
<intersection>-58 25</intersection>
<intersection>-53 21</intersection>
<intersection>-38.5 24</intersection>
<intersection>-32.5 20</intersection>
<intersection>-27 22</intersection>
<intersection>3 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>94,-69.5,95.5,-69.5</points>
<connection>
<GID>192</GID>
<name>SEL_0</name></connection>
<intersection>94 4</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>94,-82.5,94.5,-82.5</points>
<connection>
<GID>193</GID>
<name>SEL_0</name></connection>
<intersection>94 4</intersection>
<intersection>94.5 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>94.5,-99,94.5,-82.5</points>
<connection>
<GID>194</GID>
<name>SEL_0</name></connection>
<connection>
<GID>195</GID>
<name>SEL_0</name></connection>
<intersection>-99 15</intersection>
<intersection>-82.5 12</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>94.5,-99,95,-99</points>
<connection>
<GID>196</GID>
<name>SEL_0</name></connection>
<intersection>94.5 13</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>94,-32.5,94.5,-32.5</points>
<connection>
<GID>148</GID>
<name>SEL_0</name></connection>
<intersection>94 4</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>94,-53,94.5,-53</points>
<connection>
<GID>189</GID>
<name>SEL_0</name></connection>
<intersection>94 4</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>94,-27,94.5,-27</points>
<connection>
<GID>146</GID>
<name>SEL_0</name></connection>
<intersection>94 4</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>94,-38.5,95,-38.5</points>
<connection>
<GID>188</GID>
<name>SEL_0</name></connection>
<intersection>94 4</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>94,-58,95,-58</points>
<connection>
<GID>190</GID>
<name>SEL_0</name></connection>
<intersection>94 4</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>94,-63.5,95,-63.5</points>
<connection>
<GID>191</GID>
<name>SEL_0</name></connection>
<intersection>94 4</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-24.5,100,-24.5</points>
<connection>
<GID>939</GID>
<name>IN_0</name></connection>
<connection>
<GID>144</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-23.5,89,-15</points>
<intersection>-23.5 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89,-23.5,92,-23.5</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86,-15,89,-15</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-25.5,78.5,-25</points>
<intersection>-25.5 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-25.5,92,-25.5</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-25,78.5,-25</points>
<intersection>65 3</intersection>
<intersection>78.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>65,-29.5,65,-25</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>-25 2</intersection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-57,139.5,-49</points>
<connection>
<GID>947</GID>
<name>OUT_0</name></connection>
<connection>
<GID>944</GID>
<name>SEL_0</name></connection></vsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-61.5,131,-60.5</points>
<connection>
<GID>952</GID>
<name>OUT_0</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,-60.5,137.5,-60.5</points>
<connection>
<GID>944</GID>
<name>IN_0</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-58.5,131.5,-56</points>
<connection>
<GID>959</GID>
<name>OUT_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,-58.5,137.5,-58.5</points>
<connection>
<GID>944</GID>
<name>IN_1</name></connection>
<intersection>131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-60,144.5,-59.5</points>
<intersection>-60 1</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144.5,-60,148,-60</points>
<connection>
<GID>962</GID>
<name>N_in0</name></connection>
<intersection>144.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141.5,-59.5,144.5,-59.5</points>
<connection>
<GID>944</GID>
<name>OUT</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-30.5,98.5,-29.5</points>
<intersection>-30.5 1</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,-30.5,100.5,-30.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-29.5,98.5,-29.5</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65,-30.5,92.5,-30.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<connection>
<GID>57</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-28.5,89.5,-28</points>
<intersection>-28.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-28.5,92.5,-28.5</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87,-28,89.5,-28</points>
<connection>
<GID>963</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>733</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-36,98,-35</points>
<intersection>-36 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98,-36,100,-36</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-35,98,-35</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>734</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-35.5,92.5,-35.5</points>
<intersection>75 3</intersection>
<intersection>92.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75,-35.5,75,-31.5</points>
<intersection>-35.5 1</intersection>
<intersection>-31.5 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>92.5,-36,92.5,-35.5</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>65,-31.5,75,-31.5</points>
<connection>
<GID>57</GID>
<name>OUT_2</name></connection>
<intersection>75 3</intersection></hsegment></shape></wire>
<wire>
<ID>735</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-34,90.5,-33</points>
<intersection>-34 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90.5,-34,92.5,-34</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89,-33,90.5,-33</points>
<connection>
<GID>964</GID>
<name>IN_0</name></connection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>736</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-41,98.5,-40.5</points>
<intersection>-41 2</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,-40.5,100,-40.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-41,98.5,-41</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>737</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-42,65,-32.5</points>
<connection>
<GID>57</GID>
<name>OUT_3</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65,-42,93,-42</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>738</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-40,90,-39.5</points>
<intersection>-40 1</intersection>
<intersection>-39.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-40,93,-40</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-39.5,90,-39.5</points>
<connection>
<GID>965</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>743</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96.5,-55.5,102,-55.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<connection>
<GID>189</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>744</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65,-56.5,92.5,-56.5</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>65 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>65,-60.5,65,-56.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>-56.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>749</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-54.5,85.5,-53</points>
<intersection>-54.5 1</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-54.5,92.5,-54.5</points>
<connection>
<GID>189</GID>
<name>IN_1</name></connection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78.5,-53,85.5,-53</points>
<connection>
<GID>967</GID>
<name>IN_0</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>750</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97,-60.5,101.5,-60.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<connection>
<GID>190</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>751</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65,-61.5,93,-61.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<connection>
<GID>60</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>752</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-59.5,90.5,-59</points>
<intersection>-59.5 1</intersection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90.5,-59.5,93,-59.5</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>88,-59,90.5,-59</points>
<connection>
<GID>968</GID>
<name>IN_0</name></connection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>753</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-66,99,-65.5</points>
<intersection>-66 2</intersection>
<intersection>-65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-65.5,101.5,-65.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-66,99,-66</points>
<connection>
<GID>191</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>754</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-65,92,-63.5</points>
<intersection>-65 1</intersection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,-65,93,-65</points>
<connection>
<GID>191</GID>
<name>IN_1</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90,-63.5,92,-63.5</points>
<connection>
<GID>971</GID>
<name>IN_0</name></connection>
<intersection>92 0</intersection></hsegment></shape></wire>
<wire>
<ID>755</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-67,73,-62.5</points>
<intersection>-67 1</intersection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-67,93,-67</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-62.5,73,-62.5</points>
<connection>
<GID>60</GID>
<name>OUT_2</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>756</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-72,99.5,-71.5</points>
<intersection>-72 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-71.5,102,-71.5</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-72,99.5,-72</points>
<connection>
<GID>192</GID>
<name>OUT</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>757</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-73,65.5,-63.5</points>
<intersection>-73 1</intersection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-73,93.5,-73</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-63.5,65.5,-63.5</points>
<connection>
<GID>60</GID>
<name>OUT_3</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>758</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-71,92,-70</points>
<intersection>-71 1</intersection>
<intersection>-70 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,-71,93.5,-71</points>
<connection>
<GID>192</GID>
<name>IN_1</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-70,92,-70</points>
<connection>
<GID>966</GID>
<name>IN_0</name></connection>
<intersection>92 0</intersection></hsegment></shape></wire>
<wire>
<ID>759</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-85,97.5,-84.5</points>
<intersection>-85 2</intersection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-84.5,99,-84.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96,-85,97.5,-85</points>
<connection>
<GID>193</GID>
<name>OUT</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>760</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65,-86,92,-86</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>65 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>65,-89.5,65,-86</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>-86 1</intersection></vsegment></shape></wire>
<wire>
<ID>761</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-84,87.5,-83</points>
<intersection>-84 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87.5,-84,92,-84</points>
<connection>
<GID>193</GID>
<name>IN_1</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,-83,87.5,-83</points>
<connection>
<GID>973</GID>
<name>IN_0</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>762</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-89,90.5,-87.5</points>
<intersection>-89 1</intersection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90.5,-89,92.5,-89</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>88.5,-87.5,90.5,-87.5</points>
<connection>
<GID>974</GID>
<name>IN_0</name></connection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>763</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-94.5,91.5,-93.5</points>
<intersection>-94.5 3</intersection>
<intersection>-93.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>91,-93.5,91.5,-93.5</points>
<connection>
<GID>975</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>91.5,-94.5,92.5,-94.5</points>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>764</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-100.5,91,-100</points>
<intersection>-100.5 1</intersection>
<intersection>-100 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91,-100.5,93,-100.5</points>
<connection>
<GID>196</GID>
<name>IN_1</name></connection>
<intersection>91 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89,-100,91,-100</points>
<connection>
<GID>972</GID>
<name>IN_0</name></connection>
<intersection>91 0</intersection></hsegment></shape></wire>
<wire>
<ID>765</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-102.5,65.5,-92.5</points>
<intersection>-102.5 1</intersection>
<intersection>-92.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-102.5,93,-102.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-92.5,65.5,-92.5</points>
<connection>
<GID>61</GID>
<name>OUT_3</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>766</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97,-101.5,101,-101.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<connection>
<GID>196</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>767</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-96,98.5,-95.5</points>
<intersection>-96 1</intersection>
<intersection>-95.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,-96,100.5,-96</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-95.5,98.5,-95.5</points>
<connection>
<GID>195</GID>
<name>OUT</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>768</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-96.5,78.5,-91.5</points>
<intersection>-96.5 1</intersection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-96.5,92.5,-96.5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-91.5,78.5,-91.5</points>
<connection>
<GID>61</GID>
<name>OUT_2</name></connection>
<intersection>78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>769</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96.5,-90,99,-90</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<connection>
<GID>194</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>770</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-91,78.5,-90.5</points>
<intersection>-91 1</intersection>
<intersection>-90.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-91,92.5,-91</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-90.5,78.5,-90.5</points>
<connection>
<GID>61</GID>
<name>OUT_1</name></connection>
<intersection>78.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-26.8962,58.4913,395.032,-159.117</PageViewport>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>140,69.5</position>
<gparam>LABEL_TEXT Prof.  Angelo Zanini / Nuncio Perrella</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>17</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>178.5,43.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>4 </input>
<input>
<ID>IN_3</ID>5 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>169.5,39.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_IR</lparam></gate>
<gate>
<ID>19</ID>
<type>DA_FROM</type>
<position>169.5,42.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_IR</lparam></gate>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>169.5,45.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_IR</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>169.5,48.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_IR</lparam></gate>
<gate>
<ID>22</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>158,44</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>8 </input>
<input>
<ID>IN_3</ID>9 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>23</ID>
<type>DA_FROM</type>
<position>149,40</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_IR</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>149,43</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_IR</lparam></gate>
<gate>
<ID>25</ID>
<type>DA_FROM</type>
<position>149,46</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_IR</lparam></gate>
<gate>
<ID>26</ID>
<type>DA_FROM</type>
<position>149,49</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_IR</lparam></gate>
<gate>
<ID>27</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>138,44.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>24 </input>
<input>
<ID>IN_3</ID>132 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>28</ID>
<type>DA_FROM</type>
<position>129,40.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_IR</lparam></gate>
<gate>
<ID>29</ID>
<type>DA_FROM</type>
<position>129,43.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_IR</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>129,46.5</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_IR</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>143.5,58.5</position>
<gparam>LABEL_TEXT Registrador de Instrucoes - IR</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>DE_TO</type>
<position>166,31.5</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_IR</lparam></gate>
<gate>
<ID>37</ID>
<type>DE_TO</type>
<position>166,18.5</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_IR</lparam></gate>
<gate>
<ID>38</ID>
<type>DE_TO</type>
<position>167,5.5</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_IR</lparam></gate>
<gate>
<ID>39</ID>
<type>DE_TO</type>
<position>167,-7.5</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_IR</lparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>167,-20.5</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_IR</lparam></gate>
<gate>
<ID>41</ID>
<type>DE_TO</type>
<position>167,-32.5</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_IR</lparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>167,-45.5</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_IR</lparam></gate>
<gate>
<ID>43</ID>
<type>DE_TO</type>
<position>167,-58.5</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_IR</lparam></gate>
<gate>
<ID>56</ID>
<type>DE_TO</type>
<position>167.5,-71.5</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_IR</lparam></gate>
<gate>
<ID>58</ID>
<type>DE_TO</type>
<position>167,-84.5</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_IR</lparam></gate>
<gate>
<ID>59</ID>
<type>DE_TO</type>
<position>167,-97.5</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_IR</lparam></gate>
<gate>
<ID>72</ID>
<type>DE_TO</type>
<position>167.5,-111.5</position>
<input>
<ID>IN_0</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_IR</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_DFF_LOW_NT</type>
<position>159,-113.5</position>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUT_0</ID>131 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>854</ID>
<type>AA_LABEL</type>
<position>237,13</position>
<gparam>LABEL_TEXT Sinais de Controle</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>855</ID>
<type>AA_LABEL</type>
<position>217.5,3.5</position>
<gparam>LABEL_TEXT RESET</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>856</ID>
<type>AA_LABEL</type>
<position>217.5,-1.5</position>
<gparam>LABEL_TEXT WR_IR</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>DA_FROM</type>
<position>150,-111.5</position>
<input>
<ID>IN_0</ID>130 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD11</lparam></gate>
<gate>
<ID>91</ID>
<type>DA_FROM</type>
<position>129,49.5</position>
<input>
<ID>IN_0</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_IR</lparam></gate>
<gate>
<ID>874</ID>
<type>DE_TO</type>
<position>168,-126.5</position>
<input>
<ID>IN_0</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_IR</lparam></gate>
<gate>
<ID>875</ID>
<type>DE_TO</type>
<position>167.5,-139.5</position>
<input>
<ID>IN_0</ID>695 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_IR</lparam></gate>
<gate>
<ID>876</ID>
<type>DE_TO</type>
<position>167.5,-152.5</position>
<input>
<ID>IN_0</ID>699 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_IR</lparam></gate>
<gate>
<ID>877</ID>
<type>DE_TO</type>
<position>168,-166.5</position>
<input>
<ID>IN_0</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_IR</lparam></gate>
<gate>
<ID>878</ID>
<type>AE_DFF_LOW_NT</type>
<position>159.5,-168.5</position>
<input>
<ID>IN_0</ID>702 </input>
<output>
<ID>OUTINV_0</ID>707 </output>
<output>
<ID>OUT_0</ID>703 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>879</ID>
<type>DA_FROM</type>
<position>150.5,-166.5</position>
<input>
<ID>IN_0</ID>702 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD15</lparam></gate>
<gate>
<ID>880</ID>
<type>AE_DFF_LOW_NT</type>
<position>159,-128.5</position>
<input>
<ID>IN_0</ID>696 </input>
<output>
<ID>OUTINV_0</ID>704 </output>
<output>
<ID>OUT_0</ID>694 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>881</ID>
<type>AE_DFF_LOW_NT</type>
<position>159,-141.5</position>
<input>
<ID>IN_0</ID>697 </input>
<output>
<ID>OUTINV_0</ID>705 </output>
<output>
<ID>OUT_0</ID>695 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>882</ID>
<type>AE_DFF_LOW_NT</type>
<position>159,-154.5</position>
<input>
<ID>IN_0</ID>698 </input>
<output>
<ID>OUTINV_0</ID>706 </output>
<output>
<ID>OUT_0</ID>699 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>883</ID>
<type>DA_FROM</type>
<position>150,-126.5</position>
<input>
<ID>IN_0</ID>696 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD12</lparam></gate>
<gate>
<ID>884</ID>
<type>DA_FROM</type>
<position>150,-139.5</position>
<input>
<ID>IN_0</ID>697 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD13</lparam></gate>
<gate>
<ID>885</ID>
<type>DA_FROM</type>
<position>150,-152.5</position>
<input>
<ID>IN_0</ID>698 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD14</lparam></gate>
<gate>
<ID>886</ID>
<type>DE_TO</type>
<position>168,-129.5</position>
<input>
<ID>IN_0</ID>704 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D12_IR</lparam></gate>
<gate>
<ID>887</ID>
<type>DE_TO</type>
<position>167.5,-142.5</position>
<input>
<ID>IN_0</ID>705 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D13_IR</lparam></gate>
<gate>
<ID>888</ID>
<type>DE_TO</type>
<position>167.5,-155.5</position>
<input>
<ID>IN_0</ID>706 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D14_IR</lparam></gate>
<gate>
<ID>889</ID>
<type>DE_TO</type>
<position>168,-169.5</position>
<input>
<ID>IN_0</ID>707 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D15_IR</lparam></gate>
<gate>
<ID>891</ID>
<type>AA_LABEL</type>
<position>203,-149.5</position>
<gparam>LABEL_TEXT Decodifica�ao de Instrucoes</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>145.5,81</position>
<gparam>LABEL_TEXT PROCESSADOR BIP IMT - MAUA 2022</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>159</ID>
<type>AE_DFF_LOW_NT</type>
<position>158.5,29.5</position>
<input>
<ID>IN_0</ID>97 </input>
<output>
<ID>OUT_0</ID>73 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>160</ID>
<type>AE_DFF_LOW_NT</type>
<position>158.5,16.5</position>
<input>
<ID>IN_0</ID>98 </input>
<output>
<ID>OUT_0</ID>84 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>161</ID>
<type>AE_DFF_LOW_NT</type>
<position>158.5,3.5</position>
<input>
<ID>IN_0</ID>99 </input>
<output>
<ID>OUT_0</ID>85 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>162</ID>
<type>AE_DFF_LOW_NT</type>
<position>158.5,-9.5</position>
<input>
<ID>IN_0</ID>100 </input>
<output>
<ID>OUT_0</ID>90 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>163</ID>
<type>AE_DFF_LOW_NT</type>
<position>158.5,-22.5</position>
<input>
<ID>IN_0</ID>101 </input>
<output>
<ID>OUT_0</ID>91 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>164</ID>
<type>AE_DFF_LOW_NT</type>
<position>158.5,-34.5</position>
<input>
<ID>IN_0</ID>102 </input>
<output>
<ID>OUT_0</ID>92 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>165</ID>
<type>AE_DFF_LOW_NT</type>
<position>158.5,-47.5</position>
<input>
<ID>IN_0</ID>103 </input>
<output>
<ID>OUT_0</ID>93 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>166</ID>
<type>AE_DFF_LOW_NT</type>
<position>158.5,-60.5</position>
<input>
<ID>IN_0</ID>104 </input>
<output>
<ID>OUT_0</ID>94 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>167</ID>
<type>AE_DFF_LOW_NT</type>
<position>158.5,-73.5</position>
<input>
<ID>IN_0</ID>105 </input>
<output>
<ID>OUT_0</ID>95 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>168</ID>
<type>AE_DFF_LOW_NT</type>
<position>158.5,-86.5</position>
<input>
<ID>IN_0</ID>106 </input>
<output>
<ID>OUT_0</ID>96 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>169</ID>
<type>AE_DFF_LOW_NT</type>
<position>158.5,-99.5</position>
<input>
<ID>IN_0</ID>107 </input>
<output>
<ID>OUT_0</ID>108 </output>
<input>
<ID>clear</ID>110 </input>
<input>
<ID>clock</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>171</ID>
<type>DA_FROM</type>
<position>149.5,31.5</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD0</lparam></gate>
<gate>
<ID>172</ID>
<type>DA_FROM</type>
<position>149.5,18.5</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD1</lparam></gate>
<gate>
<ID>173</ID>
<type>DA_FROM</type>
<position>149.5,5.5</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD2</lparam></gate>
<gate>
<ID>174</ID>
<type>DA_FROM</type>
<position>149.5,-7.5</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD3</lparam></gate>
<gate>
<ID>175</ID>
<type>DA_FROM</type>
<position>149.5,-20.5</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD4</lparam></gate>
<gate>
<ID>176</ID>
<type>DA_FROM</type>
<position>149.5,-32.5</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD5</lparam></gate>
<gate>
<ID>177</ID>
<type>DA_FROM</type>
<position>149.5,-45.5</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD6</lparam></gate>
<gate>
<ID>178</ID>
<type>DA_FROM</type>
<position>149.5,-58.5</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD7</lparam></gate>
<gate>
<ID>179</ID>
<type>DA_FROM</type>
<position>149.5,-71.5</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD8</lparam></gate>
<gate>
<ID>180</ID>
<type>DA_FROM</type>
<position>149.5,-84.5</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD9</lparam></gate>
<gate>
<ID>181</ID>
<type>DA_FROM</type>
<position>149.5,-97.5</position>
<input>
<ID>IN_0</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD10</lparam></gate>
<gate>
<ID>954</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>113,44.5</position>
<input>
<ID>IN_0</ID>745 </input>
<input>
<ID>IN_1</ID>746 </input>
<input>
<ID>IN_2</ID>747 </input>
<input>
<ID>IN_3</ID>748 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>183</ID>
<type>DA_FROM</type>
<position>128.5,28.5</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WR_IR</lparam></gate>
<gate>
<ID>955</ID>
<type>DA_FROM</type>
<position>104,40.5</position>
<input>
<ID>IN_0</ID>745 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_IR</lparam></gate>
<gate>
<ID>184</ID>
<type>DA_FROM</type>
<position>128.5,24</position>
<input>
<ID>IN_0</ID>110 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RESET</lparam></gate>
<gate>
<ID>956</ID>
<type>DA_FROM</type>
<position>104,43.5</position>
<input>
<ID>IN_0</ID>746 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_IR</lparam></gate>
<gate>
<ID>957</ID>
<type>DA_FROM</type>
<position>104,46.5</position>
<input>
<ID>IN_0</ID>747 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_IR</lparam></gate>
<gate>
<ID>958</ID>
<type>DA_FROM</type>
<position>104,49.5</position>
<input>
<ID>IN_0</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_IR</lparam></gate>
<gate>
<ID>960</ID>
<type>AA_LABEL</type>
<position>107,37.5</position>
<gparam>LABEL_TEXT Instrucao</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173.5,39.5,173.5,42.5</points>
<intersection>39.5 2</intersection>
<intersection>42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173.5,42.5,175.5,42.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>173.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>171.5,39.5,173.5,39.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>173.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172.5,42.5,172.5,43.5</points>
<intersection>42.5 2</intersection>
<intersection>43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172.5,43.5,175.5,43.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>172.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>171.5,42.5,172.5,42.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>172.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172.5,44.5,172.5,45.5</points>
<intersection>44.5 1</intersection>
<intersection>45.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172.5,44.5,175.5,44.5</points>
<connection>
<GID>17</GID>
<name>IN_2</name></connection>
<intersection>172.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>171.5,45.5,172.5,45.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>172.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173.5,45.5,173.5,48.5</points>
<intersection>45.5 1</intersection>
<intersection>48.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173.5,45.5,175.5,45.5</points>
<connection>
<GID>17</GID>
<name>IN_3</name></connection>
<intersection>173.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>171.5,48.5,173.5,48.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>173.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,40,153,43</points>
<intersection>40 2</intersection>
<intersection>43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>153,43,155,43</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>153 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,40,153,40</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>153 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,43,152,44</points>
<intersection>43 2</intersection>
<intersection>44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152,44,155,44</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,43,152,43</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,45,152,46</points>
<intersection>45 1</intersection>
<intersection>46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152,45,155,45</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,46,152,46</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,46,153,49</points>
<intersection>46 1</intersection>
<intersection>49 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>153,46,155,46</points>
<connection>
<GID>22</GID>
<name>IN_3</name></connection>
<intersection>153 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,49,153,49</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>153 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,40.5,133,43.5</points>
<intersection>40.5 2</intersection>
<intersection>43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,43.5,135,43.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131,40.5,133,40.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,43.5,132,44.5</points>
<intersection>43.5 2</intersection>
<intersection>44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,44.5,135,44.5</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131,43.5,132,43.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,45.5,132,46.5</points>
<intersection>45.5 1</intersection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,45.5,135,45.5</points>
<connection>
<GID>27</GID>
<name>IN_2</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131,46.5,132,46.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,31.5,164,31.5</points>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,18.5,164,18.5</points>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,5.5,165,5.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,-7.5,165,-7.5</points>
<connection>
<GID>162</GID>
<name>OUT_0</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,-20.5,165,-20.5</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,-32.5,165,-32.5</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<connection>
<GID>41</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,-45.5,165,-45.5</points>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<connection>
<GID>42</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,-58.5,165,-58.5</points>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<connection>
<GID>43</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,-71.5,165.5,-71.5</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<connection>
<GID>56</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,-84.5,165,-84.5</points>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection>
<connection>
<GID>58</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,31.5,155.5,31.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<connection>
<GID>171</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,18.5,155.5,18.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<connection>
<GID>172</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,5.5,155.5,5.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<connection>
<GID>161</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,-7.5,155.5,-7.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<connection>
<GID>174</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,-20.5,155.5,-20.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<connection>
<GID>175</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,-32.5,155.5,-32.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<connection>
<GID>176</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,-45.5,155.5,-45.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<connection>
<GID>177</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,-58.5,155.5,-58.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,-71.5,155.5,-71.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<connection>
<GID>179</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,-84.5,155.5,-84.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<connection>
<GID>180</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,-97.5,155.5,-97.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<connection>
<GID>181</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,-97.5,165,-97.5</points>
<connection>
<GID>169</GID>
<name>OUT_0</name></connection>
<connection>
<GID>59</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>130.5,28.5,155.5,28.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<connection>
<GID>159</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>136.5,-169.5,136.5,28.5</points>
<intersection>-169.5 30</intersection>
<intersection>-155.5 36</intersection>
<intersection>-142.5 34</intersection>
<intersection>-129.5 32</intersection>
<intersection>-114.5 28</intersection>
<intersection>-100.5 23</intersection>
<intersection>-87.5 21</intersection>
<intersection>-74.5 19</intersection>
<intersection>-61.5 17</intersection>
<intersection>-48.5 15</intersection>
<intersection>-35.5 13</intersection>
<intersection>-23.5 11</intersection>
<intersection>-10.5 9</intersection>
<intersection>2.5 7</intersection>
<intersection>15.5 4</intersection>
<intersection>28.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>136.5,15.5,155.5,15.5</points>
<connection>
<GID>160</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>136.5,2.5,155.5,2.5</points>
<connection>
<GID>161</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>136.5,-10.5,155.5,-10.5</points>
<connection>
<GID>162</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>136.5,-23.5,155.5,-23.5</points>
<connection>
<GID>163</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>136.5,-35.5,155.5,-35.5</points>
<connection>
<GID>164</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>136.5,-48.5,155.5,-48.5</points>
<connection>
<GID>165</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>136.5,-61.5,155.5,-61.5</points>
<connection>
<GID>166</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>136.5,-74.5,155.5,-74.5</points>
<connection>
<GID>167</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>136.5,-87.5,155.5,-87.5</points>
<connection>
<GID>168</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>136.5,-100.5,155.5,-100.5</points>
<connection>
<GID>169</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>136.5,-114.5,156,-114.5</points>
<connection>
<GID>74</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>136.5,-169.5,156.5,-169.5</points>
<connection>
<GID>878</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>136.5,-129.5,156,-129.5</points>
<connection>
<GID>880</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>136.5,-142.5,156,-142.5</points>
<connection>
<GID>881</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>136.5,-155.5,156,-155.5</points>
<connection>
<GID>882</GID>
<name>clock</name></connection>
<intersection>136.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>130.5,24,158.5,24</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection>
<intersection>158.5 63</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-174,133.5,24</points>
<intersection>-174 49</intersection>
<intersection>-160 48</intersection>
<intersection>-146.5 51</intersection>
<intersection>-134 53</intersection>
<intersection>-118.5 43</intersection>
<intersection>-104.5 28</intersection>
<intersection>-91.5 26</intersection>
<intersection>-78.5 24</intersection>
<intersection>-65.5 22</intersection>
<intersection>-52.5 20</intersection>
<intersection>-39.5 18</intersection>
<intersection>-27.5 16</intersection>
<intersection>-14.5 14</intersection>
<intersection>-1.5 12</intersection>
<intersection>11 58</intersection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>133.5,-1.5,158.5,-1.5</points>
<intersection>133.5 2</intersection>
<intersection>158.5 39</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>133.5,-14.5,158.5,-14.5</points>
<intersection>133.5 2</intersection>
<intersection>158.5 38</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>133.5,-27.5,158.5,-27.5</points>
<intersection>133.5 2</intersection>
<intersection>158.5 37</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>133.5,-39.5,158.5,-39.5</points>
<intersection>133.5 2</intersection>
<intersection>158.5 36</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>133.5,-52.5,158.5,-52.5</points>
<intersection>133.5 2</intersection>
<intersection>158.5 35</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>133.5,-65.5,158.5,-65.5</points>
<intersection>133.5 2</intersection>
<intersection>158.5 34</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>133.5,-78.5,158.5,-78.5</points>
<intersection>133.5 2</intersection>
<intersection>158.5 33</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>133.5,-91.5,158.5,-91.5</points>
<intersection>133.5 2</intersection>
<intersection>158.5 32</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>133.5,-104.5,158.5,-104.5</points>
<intersection>133.5 2</intersection>
<intersection>158.5 31</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>158.5,-104.5,158.5,-103.5</points>
<connection>
<GID>169</GID>
<name>clear</name></connection>
<intersection>-104.5 28</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>158.5,-91.5,158.5,-90.5</points>
<connection>
<GID>168</GID>
<name>clear</name></connection>
<intersection>-91.5 26</intersection></vsegment>
<vsegment>
<ID>33</ID>
<points>158.5,-78.5,158.5,-77.5</points>
<connection>
<GID>167</GID>
<name>clear</name></connection>
<intersection>-78.5 24</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>158.5,-65.5,158.5,-64.5</points>
<connection>
<GID>166</GID>
<name>clear</name></connection>
<intersection>-65.5 22</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>158.5,-52.5,158.5,-51.5</points>
<connection>
<GID>165</GID>
<name>clear</name></connection>
<intersection>-52.5 20</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>158.5,-39.5,158.5,-38.5</points>
<connection>
<GID>164</GID>
<name>clear</name></connection>
<intersection>-39.5 18</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>158.5,-27.5,158.5,-26.5</points>
<connection>
<GID>163</GID>
<name>clear</name></connection>
<intersection>-27.5 16</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>158.5,-14.5,158.5,-13.5</points>
<connection>
<GID>162</GID>
<name>clear</name></connection>
<intersection>-14.5 14</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>158.5,-1.5,158.5,-0.5</points>
<connection>
<GID>161</GID>
<name>clear</name></connection>
<intersection>-1.5 12</intersection></vsegment>
<hsegment>
<ID>43</ID>
<points>133.5,-118.5,159,-118.5</points>
<intersection>133.5 2</intersection>
<intersection>159 44</intersection></hsegment>
<vsegment>
<ID>44</ID>
<points>159,-118.5,159,-117.5</points>
<connection>
<GID>74</GID>
<name>clear</name></connection>
<intersection>-118.5 43</intersection></vsegment>
<hsegment>
<ID>48</ID>
<points>133.5,-160,159,-160</points>
<intersection>133.5 2</intersection>
<intersection>159 56</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>133.5,-174,159.5,-174</points>
<intersection>133.5 2</intersection>
<intersection>159.5 57</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>133.5,-146.5,159,-146.5</points>
<intersection>133.5 2</intersection>
<intersection>159 55</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>133.5,-134,159,-134</points>
<intersection>133.5 2</intersection>
<intersection>159 54</intersection></hsegment>
<vsegment>
<ID>54</ID>
<points>159,-134,159,-132.5</points>
<connection>
<GID>880</GID>
<name>clear</name></connection>
<intersection>-134 53</intersection></vsegment>
<vsegment>
<ID>55</ID>
<points>159,-146.5,159,-145.5</points>
<connection>
<GID>881</GID>
<name>clear</name></connection>
<intersection>-146.5 51</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>159,-160,159,-158.5</points>
<connection>
<GID>882</GID>
<name>clear</name></connection>
<intersection>-160 48</intersection></vsegment>
<vsegment>
<ID>57</ID>
<points>159.5,-174,159.5,-172.5</points>
<connection>
<GID>878</GID>
<name>clear</name></connection>
<intersection>-174 49</intersection></vsegment>
<hsegment>
<ID>58</ID>
<points>133.5,11,158.5,11</points>
<intersection>133.5 2</intersection>
<intersection>158.5 64</intersection></hsegment>
<vsegment>
<ID>63</ID>
<points>158.5,24,158.5,25.5</points>
<connection>
<GID>159</GID>
<name>clear</name></connection>
<intersection>24 1</intersection></vsegment>
<vsegment>
<ID>64</ID>
<points>158.5,11,158.5,12.5</points>
<connection>
<GID>160</GID>
<name>clear</name></connection>
<intersection>11 58</intersection></vsegment></shape></wire>
<wire>
<ID>694</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-126.5,166,-126.5</points>
<connection>
<GID>880</GID>
<name>OUT_0</name></connection>
<connection>
<GID>874</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>695</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-139.5,165.5,-139.5</points>
<connection>
<GID>881</GID>
<name>OUT_0</name></connection>
<connection>
<GID>875</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>696</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>152,-126.5,156,-126.5</points>
<connection>
<GID>880</GID>
<name>IN_0</name></connection>
<connection>
<GID>883</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>697</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>152,-139.5,156,-139.5</points>
<connection>
<GID>881</GID>
<name>IN_0</name></connection>
<connection>
<GID>884</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>698</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>152,-152.5,156,-152.5</points>
<connection>
<GID>882</GID>
<name>IN_0</name></connection>
<connection>
<GID>885</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>699</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-152.5,165.5,-152.5</points>
<connection>
<GID>882</GID>
<name>OUT_0</name></connection>
<connection>
<GID>876</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>702</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>152.5,-166.5,156.5,-166.5</points>
<connection>
<GID>878</GID>
<name>IN_0</name></connection>
<connection>
<GID>879</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>703</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162.5,-166.5,166,-166.5</points>
<connection>
<GID>878</GID>
<name>OUT_0</name></connection>
<connection>
<GID>877</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>704</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-129.5,166,-129.5</points>
<connection>
<GID>880</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>886</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>705</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-142.5,165.5,-142.5</points>
<connection>
<GID>881</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>887</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>706</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-155.5,165.5,-155.5</points>
<connection>
<GID>882</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>888</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>707</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162.5,-169.5,166,-169.5</points>
<connection>
<GID>878</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>889</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>152,-111.5,156,-111.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<connection>
<GID>86</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-111.5,165.5,-111.5</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<connection>
<GID>72</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,46.5,133,49.5</points>
<intersection>46.5 2</intersection>
<intersection>49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,49.5,133,49.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>133,46.5,135,46.5</points>
<connection>
<GID>27</GID>
<name>IN_3</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>745</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,40.5,108,43.5</points>
<intersection>40.5 2</intersection>
<intersection>43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,43.5,110,43.5</points>
<connection>
<GID>954</GID>
<name>IN_0</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>106,40.5,108,40.5</points>
<connection>
<GID>955</GID>
<name>IN_0</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>746</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,43.5,107,44.5</points>
<intersection>43.5 2</intersection>
<intersection>44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,44.5,110,44.5</points>
<connection>
<GID>954</GID>
<name>IN_1</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>106,43.5,107,43.5</points>
<connection>
<GID>956</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>747</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,45.5,107,46.5</points>
<intersection>45.5 1</intersection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,45.5,110,45.5</points>
<connection>
<GID>954</GID>
<name>IN_2</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>106,46.5,107,46.5</points>
<connection>
<GID>957</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>748</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,46.5,108,49.5</points>
<intersection>46.5 2</intersection>
<intersection>49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,49.5,108,49.5</points>
<connection>
<GID>958</GID>
<name>IN_0</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108,46.5,110,46.5</points>
<connection>
<GID>954</GID>
<name>IN_3</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>142.408,-23.7558,450.338,-182.57</PageViewport>
<gate>
<ID>580</ID>
<type>GA_LED</type>
<position>307,-54.5</position>
<input>
<ID>N_in0</ID>146 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>582</ID>
<type>GA_LED</type>
<position>307,-61</position>
<input>
<ID>N_in0</ID>147 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>584</ID>
<type>GA_LED</type>
<position>307,-67</position>
<input>
<ID>N_in0</ID>148 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>586</ID>
<type>GA_LED</type>
<position>307,-73</position>
<input>
<ID>N_in0</ID>149 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>588</ID>
<type>GA_LED</type>
<position>307,-79</position>
<input>
<ID>N_in0</ID>150 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>590</ID>
<type>GA_LED</type>
<position>307,-85</position>
<input>
<ID>N_in0</ID>151 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>GA_LED</type>
<position>307.5,-97</position>
<input>
<ID>N_in0</ID>145 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>592</ID>
<type>GA_LED</type>
<position>307,-91.5</position>
<input>
<ID>N_in0</ID>152 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>206</ID>
<type>DE_TO</type>
<position>297,-128</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_ES</lparam></gate>
<gate>
<ID>207</ID>
<type>DE_TO</type>
<position>296,-57</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_ES</lparam></gate>
<gate>
<ID>208</ID>
<type>DE_TO</type>
<position>296,-63</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_ES</lparam></gate>
<gate>
<ID>209</ID>
<type>DE_TO</type>
<position>296.5,-69.5</position>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_ES</lparam></gate>
<gate>
<ID>210</ID>
<type>DE_TO</type>
<position>296.5,-76</position>
<input>
<ID>IN_0</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_ES</lparam></gate>
<gate>
<ID>211</ID>
<type>DE_TO</type>
<position>296.5,-82</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_ES</lparam></gate>
<gate>
<ID>213</ID>
<type>FF_GND</type>
<position>287,-138.5</position>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>215</ID>
<type>AA_LABEL</type>
<position>299.5,-46.5</position>
<gparam>LABEL_TEXT Extensao de Sinal</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>GA_LED</type>
<position>307.5,-103.5</position>
<input>
<ID>N_in0</ID>197 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>260</ID>
<type>GA_LED</type>
<position>307.5,-109.5</position>
<input>
<ID>N_in0</ID>198 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>274</ID>
<type>GA_LED</type>
<position>307.5,-115.5</position>
<input>
<ID>N_in0</ID>199 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>276</ID>
<type>GA_LED</type>
<position>307.5,-121.5</position>
<input>
<ID>N_in0</ID>200 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>280</ID>
<type>DE_TO</type>
<position>296.5,-99.5</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_ES</lparam></gate>
<gate>
<ID>282</ID>
<type>DE_TO</type>
<position>296.5,-105.5</position>
<input>
<ID>IN_0</ID>197 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_ES</lparam></gate>
<gate>
<ID>285</ID>
<type>DE_TO</type>
<position>297,-112</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_ES</lparam></gate>
<gate>
<ID>286</ID>
<type>DE_TO</type>
<position>297,-118.5</position>
<input>
<ID>IN_0</ID>199 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_ES</lparam></gate>
<gate>
<ID>287</ID>
<type>DE_TO</type>
<position>297,-124.5</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_ES</lparam></gate>
<gate>
<ID>288</ID>
<type>DA_FROM</type>
<position>290,-99.5</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_IR</lparam></gate>
<gate>
<ID>289</ID>
<type>DA_FROM</type>
<position>290,-105.5</position>
<input>
<ID>IN_0</ID>197 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_IR</lparam></gate>
<gate>
<ID>292</ID>
<type>DA_FROM</type>
<position>290.5,-112</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_IR</lparam></gate>
<gate>
<ID>293</ID>
<type>DA_FROM</type>
<position>290.5,-118.5</position>
<input>
<ID>IN_0</ID>199 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_IR</lparam></gate>
<gate>
<ID>294</ID>
<type>DA_FROM</type>
<position>290.5,-124.5</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_IR</lparam></gate>
<gate>
<ID>101</ID>
<type>DA_FROM</type>
<position>289.5,-57</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_IR</lparam></gate>
<gate>
<ID>103</ID>
<type>DA_FROM</type>
<position>289.5,-63</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_IR</lparam></gate>
<gate>
<ID>105</ID>
<type>DA_FROM</type>
<position>290,-69.5</position>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_IR</lparam></gate>
<gate>
<ID>107</ID>
<type>DA_FROM</type>
<position>290,-76</position>
<input>
<ID>IN_0</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_IR</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_LABEL</type>
<position>305,-38</position>
<gparam>LABEL_TEXT Prof.  Angelo Zanini / Nuncio Perrella</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>290,-82</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_IR</lparam></gate>
<gate>
<ID>127</ID>
<type>DA_FROM</type>
<position>290,-88</position>
<input>
<ID>IN_0</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_IR</lparam></gate>
<gate>
<ID>129</ID>
<type>DA_FROM</type>
<position>290,-94</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_IR</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>308.5,-28.5</position>
<gparam>LABEL_TEXT PROCESSADOR BIP IMT - MAUA 2022</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>156</ID>
<type>DE_TO</type>
<position>296.5,-88</position>
<input>
<ID>IN_0</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_ES</lparam></gate>
<gate>
<ID>157</ID>
<type>DE_TO</type>
<position>296.5,-94</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_ES</lparam></gate>
<gate>
<ID>170</ID>
<type>DE_TO</type>
<position>297,-131</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_ES</lparam></gate>
<gate>
<ID>182</ID>
<type>DE_TO</type>
<position>297.5,-134</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_ES</lparam></gate>
<gate>
<ID>185</ID>
<type>DE_TO</type>
<position>297,-137</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_ES</lparam></gate>
<wire>
<ID>197</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292,-105.5,294.5,-105.5</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>293 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>293,-105.5,293,-103.5</points>
<intersection>-105.5 1</intersection>
<intersection>-103.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>293,-103.5,306.5,-103.5</points>
<connection>
<GID>245</GID>
<name>N_in0</name></connection>
<intersection>293 8</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292.5,-112,295,-112</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>293 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>293,-112,293,-109.5</points>
<intersection>-112 1</intersection>
<intersection>-109.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>293,-109.5,306.5,-109.5</points>
<connection>
<GID>260</GID>
<name>N_in0</name></connection>
<intersection>293 6</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292.5,-118.5,295,-118.5</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>293 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>293,-118.5,293,-115.5</points>
<intersection>-118.5 1</intersection>
<intersection>-115.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>293,-115.5,306.5,-115.5</points>
<connection>
<GID>274</GID>
<name>N_in0</name></connection>
<intersection>293 10</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292.5,-124.5,295,-124.5</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>293 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>293,-124.5,293,-121.5</points>
<intersection>-124.5 1</intersection>
<intersection>-121.5 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>293,-121.5,306.5,-121.5</points>
<connection>
<GID>276</GID>
<name>N_in0</name></connection>
<intersection>293 16</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292,-99.5,294.5,-99.5</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>293 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>293,-99.5,293,-97</points>
<intersection>-99.5 1</intersection>
<intersection>-97 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>293,-97,306.5,-97</points>
<connection>
<GID>13</GID>
<name>N_in0</name></connection>
<intersection>293 2</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>291.5,-57,294,-57</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>293 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>293,-57,293,-54.5</points>
<intersection>-57 1</intersection>
<intersection>-54.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>293,-54.5,306,-54.5</points>
<connection>
<GID>580</GID>
<name>N_in0</name></connection>
<intersection>293 2</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>291.5,-63,294,-63</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>293 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>293,-63,293,-61</points>
<intersection>-63 1</intersection>
<intersection>-61 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>293,-61,306,-61</points>
<connection>
<GID>582</GID>
<name>N_in0</name></connection>
<intersection>293 8</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292,-69.5,294.5,-69.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>293 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>293,-69.5,293,-67</points>
<intersection>-69.5 1</intersection>
<intersection>-67 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>293,-67,306,-67</points>
<connection>
<GID>584</GID>
<name>N_in0</name></connection>
<intersection>293 6</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292,-76,294.5,-76</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>293 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>293,-76,293,-73</points>
<intersection>-76 1</intersection>
<intersection>-73 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>293,-73,306,-73</points>
<connection>
<GID>586</GID>
<name>N_in0</name></connection>
<intersection>293 10</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292,-82,294.5,-82</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>293 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>293,-82,293,-79</points>
<intersection>-82 1</intersection>
<intersection>-79 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>293,-79,306,-79</points>
<connection>
<GID>588</GID>
<name>N_in0</name></connection>
<intersection>293 16</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292,-88,294.5,-88</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>293 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>293,-88,293,-85</points>
<intersection>-88 1</intersection>
<intersection>-85 21</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>293,-85,306,-85</points>
<connection>
<GID>590</GID>
<name>N_in0</name></connection>
<intersection>293 20</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292,-94,294.5,-94</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>293 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>293,-94,293,-91.5</points>
<intersection>-94 1</intersection>
<intersection>-91.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>293,-91.5,306,-91.5</points>
<connection>
<GID>592</GID>
<name>N_in0</name></connection>
<intersection>293 6</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287,-137.5,287,-128</points>
<connection>
<GID>213</GID>
<name>OUT_0</name></connection>
<intersection>-137 5</intersection>
<intersection>-134 6</intersection>
<intersection>-131 7</intersection>
<intersection>-128 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287,-128,295,-128</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>287 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>287,-137,295,-137</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>287 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>287,-134,295.5,-134</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>287 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>287,-131,295,-131</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>287 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>239.487,-95.0327,591.513,-276.589</PageViewport>
<gate>
<ID>15</ID>
<type>DA_FROM</type>
<position>293.5,-213</position>
<input>
<ID>IN_0</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_ACC_OUT</lparam></gate>
<gate>
<ID>212</ID>
<type>DA_FROM</type>
<position>293.5,-169</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_ACC_OUT</lparam></gate>
<gate>
<ID>214</ID>
<type>DE_TO</type>
<position>378.5,-199</position>
<input>
<ID>IN_0</ID>169 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_RAM</lparam></gate>
<gate>
<ID>216</ID>
<type>DE_TO</type>
<position>378.5,-202</position>
<input>
<ID>IN_0</ID>170 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_RAM</lparam></gate>
<gate>
<ID>217</ID>
<type>DE_TO</type>
<position>378.5,-205</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_RAM</lparam></gate>
<gate>
<ID>218</ID>
<type>DE_TO</type>
<position>378.5,-169</position>
<input>
<ID>IN_0</ID>159 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_RAM</lparam></gate>
<gate>
<ID>219</ID>
<type>AI_RAM_12x16</type>
<position>341,-136</position>
<input>
<ID>ADDRESS_0</ID>171 </input>
<input>
<ID>ADDRESS_1</ID>172 </input>
<input>
<ID>ADDRESS_10</ID>181 </input>
<input>
<ID>ADDRESS_11</ID>182 </input>
<input>
<ID>ADDRESS_2</ID>173 </input>
<input>
<ID>ADDRESS_3</ID>174 </input>
<input>
<ID>ADDRESS_4</ID>175 </input>
<input>
<ID>ADDRESS_5</ID>176 </input>
<input>
<ID>ADDRESS_6</ID>177 </input>
<input>
<ID>ADDRESS_7</ID>178 </input>
<input>
<ID>ADDRESS_8</ID>179 </input>
<input>
<ID>ADDRESS_9</ID>180 </input>
<input>
<ID>DATA_IN_0</ID>239 </input>
<input>
<ID>DATA_IN_1</ID>240 </input>
<input>
<ID>DATA_IN_10</ID>229 </input>
<input>
<ID>DATA_IN_11</ID>228 </input>
<input>
<ID>DATA_IN_12</ID>227 </input>
<input>
<ID>DATA_IN_13</ID>226 </input>
<input>
<ID>DATA_IN_14</ID>225 </input>
<input>
<ID>DATA_IN_15</ID>224 </input>
<input>
<ID>DATA_IN_2</ID>237 </input>
<input>
<ID>DATA_IN_3</ID>236 </input>
<input>
<ID>DATA_IN_4</ID>235 </input>
<input>
<ID>DATA_IN_5</ID>234 </input>
<input>
<ID>DATA_IN_6</ID>233 </input>
<input>
<ID>DATA_IN_7</ID>232 </input>
<input>
<ID>DATA_IN_8</ID>231 </input>
<input>
<ID>DATA_IN_9</ID>230 </input>
<output>
<ID>DATA_OUT_0</ID>239 </output>
<output>
<ID>DATA_OUT_1</ID>240 </output>
<output>
<ID>DATA_OUT_10</ID>229 </output>
<output>
<ID>DATA_OUT_11</ID>228 </output>
<output>
<ID>DATA_OUT_12</ID>227 </output>
<output>
<ID>DATA_OUT_13</ID>226 </output>
<output>
<ID>DATA_OUT_14</ID>225 </output>
<output>
<ID>DATA_OUT_15</ID>224 </output>
<output>
<ID>DATA_OUT_2</ID>237 </output>
<output>
<ID>DATA_OUT_3</ID>236 </output>
<output>
<ID>DATA_OUT_4</ID>235 </output>
<output>
<ID>DATA_OUT_5</ID>234 </output>
<output>
<ID>DATA_OUT_6</ID>233 </output>
<output>
<ID>DATA_OUT_7</ID>232 </output>
<output>
<ID>DATA_OUT_8</ID>231 </output>
<output>
<ID>DATA_OUT_9</ID>230 </output>
<input>
<ID>ENABLE_0</ID>219 </input>
<input>
<ID>write_clock</ID>890 </input>
<input>
<ID>write_enable</ID>222 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:0 55857</lparam>
<lparam>Address:1 9489</lparam>
<lparam>Address:8 8</lparam>
<lparam>Address:9 9</lparam>
<lparam>Address:10 10</lparam>
<lparam>Address:11 11</lparam>
<lparam>Address:12 12</lparam>
<lparam>Address:16 1107</lparam>
<lparam>Address:32 101</lparam>
<lparam>Address:33 2</lparam>
<lparam>Address:48 17</lparam>
<lparam>Address:52 2</lparam>
<lparam>Address:64 7</lparam>
<lparam>Address:112 5</lparam>
<lparam>Address:113 2</lparam>
<lparam>Address:1107 1107</lparam></gate>
<gate>
<ID>220</ID>
<type>DE_TO</type>
<position>378.5,-172</position>
<input>
<ID>IN_0</ID>160 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_RAM</lparam></gate>
<gate>
<ID>221</ID>
<type>DA_FROM</type>
<position>293,-153.5</position>
<input>
<ID>IN_0</ID>171 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_IR</lparam></gate>
<gate>
<ID>222</ID>
<type>DA_FROM</type>
<position>293,-150.5</position>
<input>
<ID>IN_0</ID>172 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_IR</lparam></gate>
<gate>
<ID>223</ID>
<type>DA_FROM</type>
<position>293,-147.5</position>
<input>
<ID>IN_0</ID>173 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_IR</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>293.5,-210.5</position>
<input>
<ID>IN_0</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_ACC_OUT</lparam></gate>
<gate>
<ID>224</ID>
<type>DA_FROM</type>
<position>293,-144.5</position>
<input>
<ID>IN_0</ID>174 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_IR</lparam></gate>
<gate>
<ID>225</ID>
<type>DE_TO</type>
<position>378.5,-175</position>
<input>
<ID>IN_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_RAM</lparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>293.5,-208</position>
<input>
<ID>IN_0</ID>142 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_ACC_OUT</lparam></gate>
<gate>
<ID>226</ID>
<type>DA_FROM</type>
<position>293,-141.5</position>
<input>
<ID>IN_0</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_IR</lparam></gate>
<gate>
<ID>227</ID>
<type>DA_FROM</type>
<position>293,-138.5</position>
<input>
<ID>IN_0</ID>176 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_IR</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>293.5,-205</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_ACC_OUT</lparam></gate>
<gate>
<ID>228</ID>
<type>DA_FROM</type>
<position>293,-135.5</position>
<input>
<ID>IN_0</ID>177 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_IR</lparam></gate>
<gate>
<ID>229</ID>
<type>DA_FROM</type>
<position>293,-132.5</position>
<input>
<ID>IN_0</ID>178 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_IR</lparam></gate>
<gate>
<ID>230</ID>
<type>DE_TO</type>
<position>378.5,-178</position>
<input>
<ID>IN_0</ID>162 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_RAM</lparam></gate>
<gate>
<ID>231</ID>
<type>DA_FROM</type>
<position>293,-129.5</position>
<input>
<ID>IN_0</ID>179 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_IR</lparam></gate>
<gate>
<ID>232</ID>
<type>DA_FROM</type>
<position>293,-126.5</position>
<input>
<ID>IN_0</ID>180 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_IR</lparam></gate>
<gate>
<ID>233</ID>
<type>DA_FROM</type>
<position>293,-123.5</position>
<input>
<ID>IN_0</ID>181 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_IR</lparam></gate>
<gate>
<ID>234</ID>
<type>DA_FROM</type>
<position>293,-120.5</position>
<input>
<ID>IN_0</ID>182 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_IR</lparam></gate>
<gate>
<ID>235</ID>
<type>AA_LABEL</type>
<position>336,-109.5</position>
<gparam>LABEL_TEXT Memoria de Dados</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>236</ID>
<type>DE_TO</type>
<position>378.5,-181</position>
<input>
<ID>IN_0</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_RAM</lparam></gate>
<gate>
<ID>237</ID>
<type>DE_TO</type>
<position>378.5,-184</position>
<input>
<ID>IN_0</ID>164 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_RAM</lparam></gate>
<gate>
<ID>238</ID>
<type>DE_TO</type>
<position>378.5,-187</position>
<input>
<ID>IN_0</ID>165 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_RAM</lparam></gate>
<gate>
<ID>239</ID>
<type>DE_TO</type>
<position>378.5,-190</position>
<input>
<ID>IN_0</ID>166 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_RAM</lparam></gate>
<gate>
<ID>240</ID>
<type>DE_TO</type>
<position>378.5,-208</position>
<input>
<ID>IN_0</ID>184 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_RAM</lparam></gate>
<gate>
<ID>241</ID>
<type>DE_TO</type>
<position>378.5,-211</position>
<input>
<ID>IN_0</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_RAM</lparam></gate>
<gate>
<ID>242</ID>
<type>DE_TO</type>
<position>378.5,-214</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_RAM</lparam></gate>
<gate>
<ID>243</ID>
<type>DE_TO</type>
<position>378.5,-193</position>
<input>
<ID>IN_0</ID>167 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_RAM</lparam></gate>
<gate>
<ID>244</ID>
<type>DE_TO</type>
<position>378.5,-196</position>
<input>
<ID>IN_0</ID>168 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_RAM</lparam></gate>
<gate>
<ID>62</ID>
<type>DA_FROM</type>
<position>293.5,-202</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_ACC_OUT</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>293.5,-199</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_ACC_OUT</lparam></gate>
<gate>
<ID>65</ID>
<type>DA_FROM</type>
<position>293.5,-196</position>
<input>
<ID>IN_0</ID>138 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_ACC_OUT</lparam></gate>
<gate>
<ID>66</ID>
<type>DA_FROM</type>
<position>293.5,-193</position>
<input>
<ID>IN_0</ID>137 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_ACC_OUT</lparam></gate>
<gate>
<ID>259</ID>
<type>AA_LABEL</type>
<position>332,-86</position>
<gparam>LABEL_TEXT PROCESSADOR BIP IMT - MAUA 2022</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>68</ID>
<type>DA_FROM</type>
<position>293.5,-190</position>
<input>
<ID>IN_0</ID>136 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_ACC_OUT</lparam></gate>
<gate>
<ID>70</ID>
<type>DA_FROM</type>
<position>293.5,-187</position>
<input>
<ID>IN_0</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_ACC_OUT</lparam></gate>
<gate>
<ID>267</ID>
<type>DA_FROM</type>
<position>366,-129.5</position>
<input>
<ID>IN_0</ID>889 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>269</ID>
<type>EE_VDD</type>
<position>359.5,-138</position>
<output>
<ID>OUT_0</ID>219 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>275</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>355,-176</position>
<input>
<ID>ENABLE_0</ID>888 </input>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>240 </input>
<input>
<ID>IN_10</ID>229 </input>
<input>
<ID>IN_11</ID>228 </input>
<input>
<ID>IN_12</ID>227 </input>
<input>
<ID>IN_13</ID>226 </input>
<input>
<ID>IN_14</ID>225 </input>
<input>
<ID>IN_15</ID>224 </input>
<input>
<ID>IN_2</ID>237 </input>
<input>
<ID>IN_3</ID>236 </input>
<input>
<ID>IN_4</ID>235 </input>
<input>
<ID>IN_5</ID>234 </input>
<input>
<ID>IN_6</ID>233 </input>
<input>
<ID>IN_7</ID>232 </input>
<input>
<ID>IN_8</ID>231 </input>
<input>
<ID>IN_9</ID>230 </input>
<output>
<ID>OUT_0</ID>186 </output>
<output>
<ID>OUT_1</ID>185 </output>
<output>
<ID>OUT_10</ID>164 </output>
<output>
<ID>OUT_11</ID>163 </output>
<output>
<ID>OUT_12</ID>162 </output>
<output>
<ID>OUT_13</ID>161 </output>
<output>
<ID>OUT_14</ID>160 </output>
<output>
<ID>OUT_15</ID>159 </output>
<output>
<ID>OUT_2</ID>184 </output>
<output>
<ID>OUT_3</ID>183 </output>
<output>
<ID>OUT_4</ID>170 </output>
<output>
<ID>OUT_5</ID>169 </output>
<output>
<ID>OUT_6</ID>168 </output>
<output>
<ID>OUT_7</ID>167 </output>
<output>
<ID>OUT_8</ID>166 </output>
<output>
<ID>OUT_9</ID>165 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>277</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>320,-176</position>
<input>
<ID>ENABLE_0</ID>870 </input>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>143 </input>
<input>
<ID>IN_10</ID>134 </input>
<input>
<ID>IN_11</ID>133 </input>
<input>
<ID>IN_12</ID>129 </input>
<input>
<ID>IN_13</ID>128 </input>
<input>
<ID>IN_14</ID>127 </input>
<input>
<ID>IN_15</ID>71 </input>
<input>
<ID>IN_2</ID>142 </input>
<input>
<ID>IN_3</ID>141 </input>
<input>
<ID>IN_4</ID>140 </input>
<input>
<ID>IN_5</ID>139 </input>
<input>
<ID>IN_6</ID>138 </input>
<input>
<ID>IN_7</ID>137 </input>
<input>
<ID>IN_8</ID>136 </input>
<input>
<ID>IN_9</ID>135 </input>
<output>
<ID>OUT_0</ID>239 </output>
<output>
<ID>OUT_1</ID>240 </output>
<output>
<ID>OUT_10</ID>229 </output>
<output>
<ID>OUT_11</ID>228 </output>
<output>
<ID>OUT_12</ID>227 </output>
<output>
<ID>OUT_13</ID>226 </output>
<output>
<ID>OUT_14</ID>225 </output>
<output>
<ID>OUT_15</ID>224 </output>
<output>
<ID>OUT_2</ID>237 </output>
<output>
<ID>OUT_3</ID>236 </output>
<output>
<ID>OUT_4</ID>235 </output>
<output>
<ID>OUT_5</ID>234 </output>
<output>
<ID>OUT_6</ID>233 </output>
<output>
<ID>OUT_7</ID>232 </output>
<output>
<ID>OUT_8</ID>231 </output>
<output>
<ID>OUT_9</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>858</ID>
<type>AA_LABEL</type>
<position>426,-130</position>
<gparam>LABEL_TEXT Sinais de Controle</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>860</ID>
<type>AA_LABEL</type>
<position>408.5,-138.5</position>
<gparam>LABEL_TEXT WR_RAM</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>861</ID>
<type>AA_LABEL</type>
<position>406.5,-145.5</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>283</ID>
<type>DA_FROM</type>
<position>293.5,-166</position>
<input>
<ID>IN_0</ID>870 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WR_RAM</lparam></gate>
<gate>
<ID>284</ID>
<type>DA_FROM</type>
<position>366,-135.5</position>
<input>
<ID>IN_0</ID>222 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID WR_RAM</lparam></gate>
<gate>
<ID>92</ID>
<type>DA_FROM</type>
<position>293.5,-184</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_ACC_OUT</lparam></gate>
<gate>
<ID>123</ID>
<type>DA_FROM</type>
<position>293.5,-181</position>
<input>
<ID>IN_0</ID>133 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_ACC_OUT</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>331.5,-99.5</position>
<gparam>LABEL_TEXT Prof.  Angelo Zanini / Nuncio Perrella</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>293.5,-178</position>
<input>
<ID>IN_0</ID>129 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_ACC_OUT</lparam></gate>
<gate>
<ID>1109</ID>
<type>AA_INVERTER</type>
<position>326,-165.5</position>
<input>
<ID>IN_0</ID>870 </input>
<output>
<ID>OUT_0</ID>888 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1111</ID>
<type>AA_INVERTER</type>
<position>357,-129.5</position>
<input>
<ID>IN_0</ID>889 </input>
<output>
<ID>OUT_0</ID>890 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>154</ID>
<type>DA_FROM</type>
<position>293.5,-175</position>
<input>
<ID>IN_0</ID>128 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_ACC_OUT</lparam></gate>
<gate>
<ID>155</ID>
<type>DA_FROM</type>
<position>293.5,-172</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_ACC_OUT</lparam></gate>
<wire>
<ID>219</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350,-136.5,351.5,-136.5</points>
<connection>
<GID>219</GID>
<name>ENABLE_0</name></connection>
<intersection>351.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>351.5,-140.5,351.5,-136.5</points>
<intersection>-140.5 7</intersection>
<intersection>-136.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>351.5,-140.5,359.5,-140.5</points>
<intersection>351.5 6</intersection>
<intersection>359.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>359.5,-140.5,359.5,-139</points>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection>
<intersection>-140.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350,-135.5,364,-135.5</points>
<connection>
<GID>219</GID>
<name>write_enable</name></connection>
<connection>
<GID>284</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-168.5,353,-168.5</points>
<connection>
<GID>275</GID>
<name>IN_15</name></connection>
<connection>
<GID>277</GID>
<name>OUT_15</name></connection>
<intersection>333.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>333.5,-168.5,333.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_15</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_15</name></connection>
<intersection>-168.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-169.5,353,-169.5</points>
<connection>
<GID>275</GID>
<name>IN_14</name></connection>
<connection>
<GID>277</GID>
<name>OUT_14</name></connection>
<intersection>334.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>334.5,-169.5,334.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_14</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_14</name></connection>
<intersection>-169.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-170.5,353,-170.5</points>
<connection>
<GID>275</GID>
<name>IN_13</name></connection>
<connection>
<GID>277</GID>
<name>OUT_13</name></connection>
<intersection>335.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>335.5,-170.5,335.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_13</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_13</name></connection>
<intersection>-170.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-171.5,353,-171.5</points>
<connection>
<GID>275</GID>
<name>IN_12</name></connection>
<connection>
<GID>277</GID>
<name>OUT_12</name></connection>
<intersection>336.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>336.5,-171.5,336.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_12</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_12</name></connection>
<intersection>-171.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-172.5,353,-172.5</points>
<connection>
<GID>275</GID>
<name>IN_11</name></connection>
<connection>
<GID>277</GID>
<name>OUT_11</name></connection>
<intersection>337.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>337.5,-172.5,337.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_11</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_11</name></connection>
<intersection>-172.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-173.5,353,-173.5</points>
<connection>
<GID>275</GID>
<name>IN_10</name></connection>
<connection>
<GID>277</GID>
<name>OUT_10</name></connection>
<intersection>338.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>338.5,-173.5,338.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_10</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_10</name></connection>
<intersection>-173.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-174.5,353,-174.5</points>
<connection>
<GID>275</GID>
<name>IN_9</name></connection>
<connection>
<GID>277</GID>
<name>OUT_9</name></connection>
<intersection>339.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>339.5,-174.5,339.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_9</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_9</name></connection>
<intersection>-174.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-175.5,353,-175.5</points>
<connection>
<GID>275</GID>
<name>IN_8</name></connection>
<connection>
<GID>277</GID>
<name>OUT_8</name></connection>
<intersection>340.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>340.5,-175.5,340.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_8</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_8</name></connection>
<intersection>-175.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-176.5,353,-176.5</points>
<connection>
<GID>275</GID>
<name>IN_7</name></connection>
<connection>
<GID>277</GID>
<name>OUT_7</name></connection>
<intersection>341.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>341.5,-176.5,341.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_7</name></connection>
<intersection>-176.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-177.5,353,-177.5</points>
<connection>
<GID>275</GID>
<name>IN_6</name></connection>
<connection>
<GID>277</GID>
<name>OUT_6</name></connection>
<intersection>342.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>342.5,-177.5,342.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_6</name></connection>
<intersection>-177.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-178.5,353,-178.5</points>
<connection>
<GID>275</GID>
<name>IN_5</name></connection>
<connection>
<GID>277</GID>
<name>OUT_5</name></connection>
<intersection>343.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>343.5,-178.5,343.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_5</name></connection>
<intersection>-178.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-179.5,353,-179.5</points>
<connection>
<GID>275</GID>
<name>IN_4</name></connection>
<connection>
<GID>277</GID>
<name>OUT_4</name></connection>
<intersection>344.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>344.5,-179.5,344.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_4</name></connection>
<intersection>-179.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-180.5,353,-180.5</points>
<connection>
<GID>275</GID>
<name>IN_3</name></connection>
<connection>
<GID>277</GID>
<name>OUT_3</name></connection>
<intersection>345.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>345.5,-180.5,345.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_3</name></connection>
<intersection>-180.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-181.5,353,-181.5</points>
<connection>
<GID>275</GID>
<name>IN_2</name></connection>
<connection>
<GID>277</GID>
<name>OUT_2</name></connection>
<intersection>346.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>346.5,-181.5,346.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_2</name></connection>
<intersection>-181.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-183.5,353,-183.5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<connection>
<GID>277</GID>
<name>OUT_0</name></connection>
<intersection>348.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>348.5,-183.5,348.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_0</name></connection>
<intersection>-183.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>322,-182.5,353,-182.5</points>
<connection>
<GID>275</GID>
<name>IN_1</name></connection>
<connection>
<GID>277</GID>
<name>OUT_1</name></connection>
<intersection>347.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>347.5,-182.5,347.5,-147</points>
<connection>
<GID>219</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>219</GID>
<name>DATA_IN_1</name></connection>
<intersection>-182.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-169,302,-168.5</points>
<intersection>-169 2</intersection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302,-168.5,318,-168.5</points>
<connection>
<GID>277</GID>
<name>IN_15</name></connection>
<intersection>302 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295.5,-169,302,-169</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>302 0</intersection></hsegment></shape></wire>
<wire>
<ID>870</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>295.5,-165.5,323,-165.5</points>
<connection>
<GID>1109</GID>
<name>IN_0</name></connection>
<intersection>295.5 12</intersection>
<intersection>320 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>320,-167,320,-165.5</points>
<connection>
<GID>277</GID>
<name>ENABLE_0</name></connection>
<intersection>-165.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>295.5,-166,295.5,-165.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>-165.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>888</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,-167,355,-165.5</points>
<connection>
<GID>275</GID>
<name>ENABLE_0</name></connection>
<intersection>-165.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>329,-165.5,355,-165.5</points>
<connection>
<GID>1109</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment></shape></wire>
<wire>
<ID>889</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>360,-129.5,364,-129.5</points>
<connection>
<GID>1111</GID>
<name>IN_0</name></connection>
<connection>
<GID>267</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>890</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351.5,-134.5,351.5,-129.5</points>
<intersection>-134.5 1</intersection>
<intersection>-129.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350,-134.5,351.5,-134.5</points>
<connection>
<GID>219</GID>
<name>write_clock</name></connection>
<intersection>351.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351.5,-129.5,354,-129.5</points>
<connection>
<GID>1111</GID>
<name>OUT_0</name></connection>
<intersection>351.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303,-172,303,-169.5</points>
<intersection>-172 2</intersection>
<intersection>-169.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303,-169.5,318,-169.5</points>
<connection>
<GID>277</GID>
<name>IN_14</name></connection>
<intersection>303 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295.5,-172,303,-172</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>303 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,-175,304,-170.5</points>
<intersection>-175 2</intersection>
<intersection>-170.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-170.5,318,-170.5</points>
<connection>
<GID>277</GID>
<name>IN_13</name></connection>
<intersection>304 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295.5,-175,304,-175</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>305,-178,305,-171.5</points>
<intersection>-178 1</intersection>
<intersection>-171.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-178,305,-178</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>305 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>305,-171.5,318,-171.5</points>
<connection>
<GID>277</GID>
<name>IN_12</name></connection>
<intersection>305 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>306,-181,306,-172.5</points>
<intersection>-181 1</intersection>
<intersection>-172.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-181,306,-181</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>306 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>306,-172.5,318,-172.5</points>
<connection>
<GID>277</GID>
<name>IN_11</name></connection>
<intersection>306 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307,-184,307,-173.5</points>
<intersection>-184 1</intersection>
<intersection>-173.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-184,307,-184</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>307 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>307,-173.5,318,-173.5</points>
<connection>
<GID>277</GID>
<name>IN_10</name></connection>
<intersection>307 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308,-187,308,-174.5</points>
<intersection>-187 1</intersection>
<intersection>-174.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-187,308,-187</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308,-174.5,318,-174.5</points>
<connection>
<GID>277</GID>
<name>IN_9</name></connection>
<intersection>308 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-190,309,-175.5</points>
<intersection>-190 1</intersection>
<intersection>-175.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-190,309,-190</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>309 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309,-175.5,318,-175.5</points>
<connection>
<GID>277</GID>
<name>IN_8</name></connection>
<intersection>309 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,-193,310,-176.5</points>
<intersection>-193 1</intersection>
<intersection>-176.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-193,310,-193</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>310,-176.5,318,-176.5</points>
<connection>
<GID>277</GID>
<name>IN_7</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-196,311,-177.5</points>
<intersection>-196 1</intersection>
<intersection>-177.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-196,311,-196</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>311 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>311,-177.5,318,-177.5</points>
<connection>
<GID>277</GID>
<name>IN_6</name></connection>
<intersection>311 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312,-199,312,-178.5</points>
<intersection>-199 1</intersection>
<intersection>-178.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-199,312,-199</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>312 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>312,-178.5,318,-178.5</points>
<connection>
<GID>277</GID>
<name>IN_5</name></connection>
<intersection>312 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313,-202,313,-179.5</points>
<intersection>-202 1</intersection>
<intersection>-179.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-202,313,-202</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>313 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>313,-179.5,318,-179.5</points>
<connection>
<GID>277</GID>
<name>IN_4</name></connection>
<intersection>313 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314,-205,314,-180.5</points>
<intersection>-205 2</intersection>
<intersection>-180.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,-180.5,318,-180.5</points>
<connection>
<GID>277</GID>
<name>IN_3</name></connection>
<intersection>314 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295.5,-205,314,-205</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>314 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>315,-208,315,-181.5</points>
<intersection>-208 1</intersection>
<intersection>-181.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-208,315,-208</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>315 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>315,-181.5,318,-181.5</points>
<connection>
<GID>277</GID>
<name>IN_2</name></connection>
<intersection>315 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316,-210.5,316,-182.5</points>
<intersection>-210.5 1</intersection>
<intersection>-182.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-210.5,316,-210.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>316 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>316,-182.5,318,-182.5</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>316 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317,-213,317,-183.5</points>
<intersection>-213 1</intersection>
<intersection>-183.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-213,317,-213</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>317 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>317,-183.5,318,-183.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>317 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>357,-168.5,373,-168.5</points>
<connection>
<GID>275</GID>
<name>OUT_15</name></connection>
<intersection>373 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>373,-169,373,-168.5</points>
<intersection>-169 4</intersection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>373,-169,376.5,-169</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>373 3</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-172,372,-169.5</points>
<intersection>-172 1</intersection>
<intersection>-169.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>372,-172,376.5,-172</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-169.5,372,-169.5</points>
<connection>
<GID>275</GID>
<name>OUT_14</name></connection>
<intersection>372 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>371,-175,371,-170.5</points>
<intersection>-175 1</intersection>
<intersection>-170.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>371,-175,376.5,-175</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>371 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-170.5,371,-170.5</points>
<connection>
<GID>275</GID>
<name>OUT_13</name></connection>
<intersection>371 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>370,-178,370,-171.5</points>
<intersection>-178 1</intersection>
<intersection>-171.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>370,-178,376.5,-178</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>370 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-171.5,370,-171.5</points>
<connection>
<GID>275</GID>
<name>OUT_12</name></connection>
<intersection>370 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369,-181,369,-172.5</points>
<intersection>-181 1</intersection>
<intersection>-172.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>369,-181,376.5,-181</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-172.5,369,-172.5</points>
<connection>
<GID>275</GID>
<name>OUT_11</name></connection>
<intersection>369 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>368,-184,368,-173.5</points>
<intersection>-184 1</intersection>
<intersection>-173.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>368,-184,376.5,-184</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>368 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-173.5,368,-173.5</points>
<connection>
<GID>275</GID>
<name>OUT_10</name></connection>
<intersection>368 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>367,-187,367,-174.5</points>
<intersection>-187 1</intersection>
<intersection>-174.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>367,-187,376.5,-187</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>367 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-174.5,367,-174.5</points>
<connection>
<GID>275</GID>
<name>OUT_9</name></connection>
<intersection>367 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366,-190,366,-175.5</points>
<intersection>-190 1</intersection>
<intersection>-175.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>366,-190,376.5,-190</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>366 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-175.5,366,-175.5</points>
<connection>
<GID>275</GID>
<name>OUT_8</name></connection>
<intersection>366 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>365,-193,365,-176.5</points>
<intersection>-193 1</intersection>
<intersection>-176.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>365,-193,376.5,-193</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>365 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-176.5,365,-176.5</points>
<connection>
<GID>275</GID>
<name>OUT_7</name></connection>
<intersection>365 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>364,-196,364,-177.5</points>
<intersection>-196 1</intersection>
<intersection>-177.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>364,-196,376.5,-196</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>364 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-177.5,364,-177.5</points>
<connection>
<GID>275</GID>
<name>OUT_6</name></connection>
<intersection>364 0</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363,-199,363,-178.5</points>
<intersection>-199 1</intersection>
<intersection>-178.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>363,-199,376.5,-199</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>363 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-178.5,363,-178.5</points>
<connection>
<GID>275</GID>
<name>OUT_5</name></connection>
<intersection>363 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>362,-202,362,-179.5</points>
<intersection>-202 1</intersection>
<intersection>-179.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>362,-202,376.5,-202</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>362 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-179.5,362,-179.5</points>
<connection>
<GID>275</GID>
<name>OUT_4</name></connection>
<intersection>362 0</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>322,-153.5,322,-141.5</points>
<intersection>-153.5 2</intersection>
<intersection>-141.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322,-141.5,332,-141.5</points>
<connection>
<GID>219</GID>
<name>ADDRESS_0</name></connection>
<intersection>322 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295,-153.5,322,-153.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>322 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321,-150.5,321,-140.5</points>
<intersection>-150.5 2</intersection>
<intersection>-140.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321,-140.5,332,-140.5</points>
<connection>
<GID>219</GID>
<name>ADDRESS_1</name></connection>
<intersection>321 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295,-150.5,321,-150.5</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>321 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320,-147.5,320,-139.5</points>
<intersection>-147.5 2</intersection>
<intersection>-139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320,-139.5,332,-139.5</points>
<connection>
<GID>219</GID>
<name>ADDRESS_2</name></connection>
<intersection>320 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295,-147.5,320,-147.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>320 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>319,-138.5,332,-138.5</points>
<connection>
<GID>219</GID>
<name>ADDRESS_3</name></connection>
<intersection>319 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>319,-144.5,319,-138.5</points>
<intersection>-144.5 7</intersection>
<intersection>-138.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>295,-144.5,319,-144.5</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>319 6</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>315.5,-137.5,332,-137.5</points>
<connection>
<GID>219</GID>
<name>ADDRESS_4</name></connection>
<intersection>315.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>315.5,-141.5,315.5,-137.5</points>
<intersection>-141.5 4</intersection>
<intersection>-137.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>295,-141.5,315.5,-141.5</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>315.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>313,-136.5,332,-136.5</points>
<connection>
<GID>219</GID>
<name>ADDRESS_5</name></connection>
<intersection>313 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>313,-138.5,313,-136.5</points>
<intersection>-138.5 4</intersection>
<intersection>-136.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>295,-138.5,313,-138.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>313 3</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>295,-135.5,332,-135.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<connection>
<GID>219</GID>
<name>ADDRESS_6</name></connection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>323,-134.5,332,-134.5</points>
<connection>
<GID>219</GID>
<name>ADDRESS_7</name></connection>
<intersection>323 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>323,-134.5,323,-132.5</points>
<intersection>-134.5 1</intersection>
<intersection>-132.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>295,-132.5,323,-132.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>323 3</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>324.5,-133.5,332,-133.5</points>
<connection>
<GID>219</GID>
<name>ADDRESS_8</name></connection>
<intersection>324.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>324.5,-133.5,324.5,-129.5</points>
<intersection>-133.5 1</intersection>
<intersection>-129.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>295,-129.5,324.5,-129.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>324.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326,-132.5,326,-126.5</points>
<intersection>-132.5 1</intersection>
<intersection>-126.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>326,-132.5,332,-132.5</points>
<connection>
<GID>219</GID>
<name>ADDRESS_9</name></connection>
<intersection>326 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295,-126.5,326,-126.5</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>326 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327,-131.5,327,-123.5</points>
<intersection>-131.5 1</intersection>
<intersection>-123.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>327,-131.5,332,-131.5</points>
<connection>
<GID>219</GID>
<name>ADDRESS_10</name></connection>
<intersection>327 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295,-123.5,327,-123.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>327 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>328,-130.5,328,-120.5</points>
<intersection>-130.5 5</intersection>
<intersection>-120.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>295,-120.5,328,-120.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>328 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>328,-130.5,332,-130.5</points>
<connection>
<GID>219</GID>
<name>ADDRESS_11</name></connection>
<intersection>328 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361,-205,361,-180.5</points>
<intersection>-205 1</intersection>
<intersection>-180.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361,-205,376.5,-205</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>361 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-180.5,361,-180.5</points>
<connection>
<GID>275</GID>
<name>OUT_3</name></connection>
<intersection>361 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>360,-208,360,-181.5</points>
<intersection>-208 1</intersection>
<intersection>-181.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360,-208,376.5,-208</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>360 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-181.5,360,-181.5</points>
<connection>
<GID>275</GID>
<name>OUT_2</name></connection>
<intersection>360 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>359,-211,359,-182.5</points>
<intersection>-211 1</intersection>
<intersection>-182.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,-211,376.5,-211</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>359 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-182.5,359,-182.5</points>
<connection>
<GID>275</GID>
<name>OUT_1</name></connection>
<intersection>359 0</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>358,-214,358,-183.5</points>
<intersection>-214 2</intersection>
<intersection>-183.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>358,-214,376.5,-214</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>358 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>357,-183.5,358,-183.5</points>
<connection>
<GID>275</GID>
<name>OUT_0</name></connection>
<intersection>358 0</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>107.422,38.4642,644.445,-238.504</PageViewport>
<gate>
<ID>389</ID>
<type>DA_FROM</type>
<position>180.5,-197.5</position>
<input>
<ID>IN_0</ID>322 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_RAM</lparam></gate>
<gate>
<ID>390</ID>
<type>DA_FROM</type>
<position>171,-195.5</position>
<input>
<ID>IN_0</ID>323 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_ES</lparam></gate>
<gate>
<ID>391</ID>
<type>DA_FROM</type>
<position>162.5,-193.5</position>
<input>
<ID>IN_0</ID>324 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_ULA</lparam></gate>
<gate>
<ID>392</ID>
<type>AE_MUX_4x1</type>
<position>233.5,-208.5</position>
<input>
<ID>IN_0</ID>328 </input>
<input>
<ID>IN_1</ID>329 </input>
<input>
<ID>IN_2</ID>330 </input>
<output>
<ID>OUT</ID>331 </output>
<input>
<ID>SEL_0</ID>327 </input>
<input>
<ID>SEL_1</ID>326 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>393</ID>
<type>DA_FROM</type>
<position>212.5,-202.5</position>
<input>
<ID>IN_0</ID>326 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>394</ID>
<type>DA_FROM</type>
<position>212.5,-199.5</position>
<input>
<ID>IN_0</ID>327 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>395</ID>
<type>DA_FROM</type>
<position>227,-211.5</position>
<input>
<ID>IN_0</ID>328 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_RAM</lparam></gate>
<gate>
<ID>396</ID>
<type>DA_FROM</type>
<position>216,-209.5</position>
<input>
<ID>IN_0</ID>329 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_ES</lparam></gate>
<gate>
<ID>397</ID>
<type>DA_FROM</type>
<position>207.5,-207.5</position>
<input>
<ID>IN_0</ID>330 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_ULA</lparam></gate>
<gate>
<ID>398</ID>
<type>AE_MUX_4x1</type>
<position>189,-221.5</position>
<input>
<ID>IN_0</ID>334 </input>
<input>
<ID>IN_1</ID>335 </input>
<input>
<ID>IN_2</ID>336 </input>
<output>
<ID>OUT</ID>337 </output>
<input>
<ID>SEL_0</ID>333 </input>
<input>
<ID>SEL_1</ID>332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>399</ID>
<type>DA_FROM</type>
<position>168,-215.5</position>
<input>
<ID>IN_0</ID>332 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>400</ID>
<type>DA_FROM</type>
<position>168,-212.5</position>
<input>
<ID>IN_0</ID>333 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>401</ID>
<type>DA_FROM</type>
<position>182.5,-224.5</position>
<input>
<ID>IN_0</ID>334 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_RAM</lparam></gate>
<gate>
<ID>402</ID>
<type>DA_FROM</type>
<position>171.5,-222.5</position>
<input>
<ID>IN_0</ID>335 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_ES</lparam></gate>
<gate>
<ID>403</ID>
<type>DA_FROM</type>
<position>163,-220.5</position>
<input>
<ID>IN_0</ID>336 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_ULA</lparam></gate>
<gate>
<ID>404</ID>
<type>AE_MUX_4x1</type>
<position>237,-234.5</position>
<input>
<ID>IN_0</ID>340 </input>
<input>
<ID>IN_1</ID>341 </input>
<input>
<ID>IN_2</ID>342 </input>
<output>
<ID>OUT</ID>343 </output>
<input>
<ID>SEL_0</ID>339 </input>
<input>
<ID>SEL_1</ID>338 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>405</ID>
<type>DA_FROM</type>
<position>215,-228.5</position>
<input>
<ID>IN_0</ID>338 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>406</ID>
<type>DA_FROM</type>
<position>215,-225.5</position>
<input>
<ID>IN_0</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>407</ID>
<type>DA_FROM</type>
<position>229.5,-237.5</position>
<input>
<ID>IN_0</ID>340 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_RAM</lparam></gate>
<gate>
<ID>1186</ID>
<type>AF_DFF_LOW</type>
<position>299,-53.5</position>
<input>
<ID>IN_0</ID>350 </input>
<output>
<ID>OUT_0</ID>953 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>954 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>408</ID>
<type>DA_FROM</type>
<position>218.5,-235.5</position>
<input>
<ID>IN_0</ID>341 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_ES</lparam></gate>
<gate>
<ID>1187</ID>
<type>DA_FROM</type>
<position>289.5,-53.5</position>
<input>
<ID>IN_0</ID>954 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>409</ID>
<type>DA_FROM</type>
<position>210,-233.5</position>
<input>
<ID>IN_0</ID>342 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_ULA</lparam></gate>
<gate>
<ID>410</ID>
<type>AE_MUX_4x1</type>
<position>189.5,-248.5</position>
<input>
<ID>IN_0</ID>346 </input>
<input>
<ID>IN_1</ID>347 </input>
<input>
<ID>IN_2</ID>348 </input>
<output>
<ID>OUT</ID>349 </output>
<input>
<ID>SEL_0</ID>345 </input>
<input>
<ID>SEL_1</ID>344 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1189</ID>
<type>DA_FROM</type>
<position>290,-65.5</position>
<input>
<ID>IN_0</ID>955 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>411</ID>
<type>DA_FROM</type>
<position>169,-242.5</position>
<input>
<ID>IN_0</ID>344 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>1190</ID>
<type>AF_DFF_LOW</type>
<position>299.5,-65.5</position>
<input>
<ID>IN_0</ID>265 </input>
<output>
<ID>OUT_0</ID>956 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>955 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>412</ID>
<type>DA_FROM</type>
<position>169,-239.5</position>
<input>
<ID>IN_0</ID>345 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>1191</ID>
<type>DA_FROM</type>
<position>288,-78</position>
<input>
<ID>IN_0</ID>957 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>413</ID>
<type>DA_FROM</type>
<position>183.5,-251.5</position>
<input>
<ID>IN_0</ID>346 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_RAM</lparam></gate>
<gate>
<ID>1192</ID>
<type>AF_DFF_LOW</type>
<position>297.5,-78</position>
<input>
<ID>IN_0</ID>271 </input>
<output>
<ID>OUT_0</ID>958 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>957 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>414</ID>
<type>DA_FROM</type>
<position>172.5,-249.5</position>
<input>
<ID>IN_0</ID>347 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_ES</lparam></gate>
<gate>
<ID>1193</ID>
<type>DA_FROM</type>
<position>288.5,-91</position>
<input>
<ID>IN_0</ID>959 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>415</ID>
<type>DA_FROM</type>
<position>164,-247.5</position>
<input>
<ID>IN_0</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_ULA</lparam></gate>
<gate>
<ID>1194</ID>
<type>AF_DFF_LOW</type>
<position>297.5,-91.5</position>
<input>
<ID>IN_0</ID>277 </input>
<output>
<ID>OUT_0</ID>960 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>959 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1195</ID>
<type>DA_FROM</type>
<position>288.5,-103.5</position>
<input>
<ID>IN_0</ID>961 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>1196</ID>
<type>AF_DFF_LOW</type>
<position>298,-103.5</position>
<input>
<ID>IN_0</ID>283 </input>
<output>
<ID>OUT_0</ID>962 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>961 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1197</ID>
<type>DA_FROM</type>
<position>288,-115.5</position>
<input>
<ID>IN_0</ID>963 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>1198</ID>
<type>AF_DFF_LOW</type>
<position>297.5,-115.5</position>
<input>
<ID>IN_0</ID>289 </input>
<output>
<ID>OUT_0</ID>964 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>963 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>420</ID>
<type>AA_LABEL</type>
<position>82,-36</position>
<gparam>LABEL_TEXT Acumulador OUT</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>1199</ID>
<type>DA_FROM</type>
<position>288,-128</position>
<input>
<ID>IN_0</ID>965 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>1200</ID>
<type>AF_DFF_LOW</type>
<position>297.5,-128</position>
<input>
<ID>IN_0</ID>295 </input>
<output>
<ID>OUT_0</ID>966 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>965 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>422</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>93,-64</position>
<input>
<ID>IN_0</ID>360 </input>
<input>
<ID>IN_1</ID>361 </input>
<input>
<ID>IN_2</ID>362 </input>
<input>
<ID>IN_3</ID>363 </input>
<input>
<ID>IN_4</ID>359 </input>
<input>
<ID>IN_5</ID>358 </input>
<input>
<ID>IN_6</ID>357 </input>
<input>
<ID>IN_7</ID>356 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 83</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1201</ID>
<type>DA_FROM</type>
<position>288.5,-142</position>
<input>
<ID>IN_0</ID>967 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>1202</ID>
<type>AF_DFF_LOW</type>
<position>298,-142</position>
<input>
<ID>IN_0</ID>301 </input>
<output>
<ID>OUT_0</ID>968 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>967 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>424</ID>
<type>DA_FROM</type>
<position>86.5,-55.5</position>
<input>
<ID>IN_0</ID>356 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D7_ACC_OUT</lparam></gate>
<gate>
<ID>1203</ID>
<type>DA_FROM</type>
<position>288.5,-155</position>
<input>
<ID>IN_0</ID>969 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>1204</ID>
<type>AF_DFF_LOW</type>
<position>298,-155</position>
<input>
<ID>IN_0</ID>307 </input>
<output>
<ID>OUT_0</ID>970 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>969 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>426</ID>
<type>DA_FROM</type>
<position>86.5,-52.5</position>
<input>
<ID>IN_0</ID>357 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D6_ACC_OUT</lparam></gate>
<gate>
<ID>1205</ID>
<type>DA_FROM</type>
<position>288.5,-167.5</position>
<input>
<ID>IN_0</ID>971 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>1206</ID>
<type>AF_DFF_LOW</type>
<position>298,-167.5</position>
<input>
<ID>IN_0</ID>313 </input>
<output>
<ID>OUT_0</ID>972 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>971 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>428</ID>
<type>DA_FROM</type>
<position>86.5,-49.5</position>
<input>
<ID>IN_0</ID>358 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D5_ACC_OUT</lparam></gate>
<gate>
<ID>1207</ID>
<type>DA_FROM</type>
<position>288,-181.5</position>
<input>
<ID>IN_0</ID>973 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>1208</ID>
<type>AF_DFF_LOW</type>
<position>297.5,-181.5</position>
<input>
<ID>IN_0</ID>319 </input>
<output>
<ID>OUT_0</ID>974 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>973 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>430</ID>
<type>DA_FROM</type>
<position>86.5,-46.5</position>
<input>
<ID>IN_0</ID>359 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D4_ACC_OUT</lparam></gate>
<gate>
<ID>1209</ID>
<type>DA_FROM</type>
<position>288.5,-195.5</position>
<input>
<ID>IN_0</ID>975 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>431</ID>
<type>DA_FROM</type>
<position>86.5,-80.5</position>
<input>
<ID>IN_0</ID>363 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D3_ACC_OUT</lparam></gate>
<gate>
<ID>1210</ID>
<type>AF_DFF_LOW</type>
<position>297.5,-195.5</position>
<input>
<ID>IN_0</ID>325 </input>
<output>
<ID>OUT_0</ID>976 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>975 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>432</ID>
<type>DA_FROM</type>
<position>86.5,-77.5</position>
<input>
<ID>IN_0</ID>362 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D2_ACC_OUT</lparam></gate>
<gate>
<ID>1211</ID>
<type>DA_FROM</type>
<position>287.5,-208.5</position>
<input>
<ID>IN_0</ID>977 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>433</ID>
<type>DA_FROM</type>
<position>86.5,-74.5</position>
<input>
<ID>IN_0</ID>361 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D1_ACC_OUT</lparam></gate>
<gate>
<ID>1212</ID>
<type>AF_DFF_LOW</type>
<position>297,-208.5</position>
<input>
<ID>IN_0</ID>331 </input>
<output>
<ID>OUT_0</ID>978 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>977 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>434</ID>
<type>DA_FROM</type>
<position>86.5,-71.5</position>
<input>
<ID>IN_0</ID>360 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D0_ACC_OUT</lparam></gate>
<gate>
<ID>1213</ID>
<type>DA_FROM</type>
<position>288,-221</position>
<input>
<ID>IN_0</ID>979 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>1214</ID>
<type>AF_DFF_LOW</type>
<position>297,-221</position>
<input>
<ID>IN_0</ID>337 </input>
<output>
<ID>OUT_0</ID>980 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>979 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1215</ID>
<type>DA_FROM</type>
<position>287.5,-235</position>
<input>
<ID>IN_0</ID>981 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>1216</ID>
<type>AF_DFF_LOW</type>
<position>297,-235</position>
<input>
<ID>IN_0</ID>343 </input>
<output>
<ID>OUT_0</ID>982 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>981 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1217</ID>
<type>DA_FROM</type>
<position>288,-249</position>
<input>
<ID>IN_0</ID>983 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>1218</ID>
<type>AF_DFF_LOW</type>
<position>297.5,-249</position>
<input>
<ID>IN_0</ID>349 </input>
<output>
<ID>OUT_0</ID>984 </output>
<input>
<ID>clear</ID>210 </input>
<input>
<ID>clock</ID>983 </input>
<input>
<ID>clock_enable</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>444</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>72,-64</position>
<input>
<ID>IN_0</ID>376 </input>
<input>
<ID>IN_1</ID>377 </input>
<input>
<ID>IN_2</ID>378 </input>
<input>
<ID>IN_3</ID>379 </input>
<input>
<ID>IN_4</ID>375 </input>
<input>
<ID>IN_5</ID>374 </input>
<input>
<ID>IN_6</ID>373 </input>
<input>
<ID>IN_7</ID>372 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>445</ID>
<type>DA_FROM</type>
<position>65.5,-55.5</position>
<input>
<ID>IN_0</ID>372 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D15_ACC_OUT</lparam></gate>
<gate>
<ID>446</ID>
<type>DA_FROM</type>
<position>65.5,-52.5</position>
<input>
<ID>IN_0</ID>373 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D14_ACC_OUT</lparam></gate>
<gate>
<ID>447</ID>
<type>DA_FROM</type>
<position>65.5,-49.5</position>
<input>
<ID>IN_0</ID>374 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D13_ACC_OUT</lparam></gate>
<gate>
<ID>448</ID>
<type>DA_FROM</type>
<position>65.5,-46.5</position>
<input>
<ID>IN_0</ID>375 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D12_ACC_OUT</lparam></gate>
<gate>
<ID>449</ID>
<type>DA_FROM</type>
<position>65.5,-80.5</position>
<input>
<ID>IN_0</ID>379 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D11_ACC_OUT</lparam></gate>
<gate>
<ID>450</ID>
<type>DA_FROM</type>
<position>65.5,-77.5</position>
<input>
<ID>IN_0</ID>378 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D10_ACC_OUT</lparam></gate>
<gate>
<ID>451</ID>
<type>DA_FROM</type>
<position>65.5,-74.5</position>
<input>
<ID>IN_0</ID>377 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D9_ACC_OUT</lparam></gate>
<gate>
<ID>452</ID>
<type>DA_FROM</type>
<position>65.5,-71.5</position>
<input>
<ID>IN_0</ID>376 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D8_ACC_OUT</lparam></gate>
<gate>
<ID>862</ID>
<type>AA_LABEL</type>
<position>80.5,-99.5</position>
<gparam>LABEL_TEXT Sinais de Controle</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>863</ID>
<type>AA_LABEL</type>
<position>65,-108.5</position>
<gparam>LABEL_TEXT SelAccSrc_0</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>866</ID>
<type>AA_LABEL</type>
<position>65,-115</position>
<gparam>LABEL_TEXT SelAccSrc_1</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>AA_LABEL</type>
<position>61,-121.5</position>
<gparam>LABEL_TEXT WR_ACC</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>AA_LABEL</type>
<position>60,-129.5</position>
<gparam>LABEL_TEXT RESET</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>205.5,-3.5</position>
<gparam>LABEL_TEXT Prof.  Angelo Zanini / Nuncio Perrella</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>204</ID>
<type>DA_FROM</type>
<position>270.5,-51.5</position>
<input>
<ID>IN_0</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WR_ACC</lparam></gate>
<gate>
<ID>1024</ID>
<type>DE_TO</type>
<position>250,-46.5</position>
<input>
<ID>IN_0</ID>350 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_ACC_IN</lparam></gate>
<gate>
<ID>246</ID>
<type>AE_MUX_4x1</type>
<position>229,-51.5</position>
<input>
<ID>IN_0</ID>257 </input>
<input>
<ID>IN_1</ID>258 </input>
<input>
<ID>IN_2</ID>259 </input>
<output>
<ID>OUT</ID>350 </output>
<input>
<ID>SEL_0</ID>256 </input>
<input>
<ID>SEL_1</ID>255 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1025</ID>
<type>DE_TO</type>
<position>241.5,-59</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_ACC_IN</lparam></gate>
<gate>
<ID>247</ID>
<type>DE_TO</type>
<position>308,-51.5</position>
<input>
<ID>IN_0</ID>953 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_ACC_OUT</lparam></gate>
<gate>
<ID>1026</ID>
<type>DE_TO</type>
<position>251.5,-71</position>
<input>
<ID>IN_0</ID>271 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_ACC_IN</lparam></gate>
<gate>
<ID>248</ID>
<type>DE_TO</type>
<position>308,-64.5</position>
<input>
<ID>IN_0</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_ACC_OUT</lparam></gate>
<gate>
<ID>1027</ID>
<type>DE_TO</type>
<position>251,-84</position>
<input>
<ID>IN_0</ID>277 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_ACC_IN</lparam></gate>
<gate>
<ID>249</ID>
<type>DE_TO</type>
<position>309,-77.5</position>
<input>
<ID>IN_0</ID>958 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_ACC_OUT</lparam></gate>
<gate>
<ID>250</ID>
<type>DE_TO</type>
<position>309,-90.5</position>
<input>
<ID>IN_0</ID>960 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_ACC_OUT</lparam></gate>
<gate>
<ID>251</ID>
<type>DE_TO</type>
<position>309,-103.5</position>
<input>
<ID>IN_0</ID>962 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_ACC_OUT</lparam></gate>
<gate>
<ID>252</ID>
<type>DE_TO</type>
<position>309,-115.5</position>
<input>
<ID>IN_0</ID>964 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_ACC_OUT</lparam></gate>
<gate>
<ID>253</ID>
<type>DE_TO</type>
<position>309,-128.5</position>
<input>
<ID>IN_0</ID>966 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_ACC_OUT</lparam></gate>
<gate>
<ID>254</ID>
<type>DE_TO</type>
<position>309,-141.5</position>
<input>
<ID>IN_0</ID>968 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_ACC_OUT</lparam></gate>
<gate>
<ID>255</ID>
<type>DE_TO</type>
<position>309.5,-154.5</position>
<input>
<ID>IN_0</ID>970 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_ACC_OUT</lparam></gate>
<gate>
<ID>256</ID>
<type>DE_TO</type>
<position>309.5,-167.5</position>
<input>
<ID>IN_0</ID>972 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_ACC_OUT</lparam></gate>
<gate>
<ID>257</ID>
<type>DE_TO</type>
<position>309,-180.5</position>
<input>
<ID>IN_0</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_ACC_OUT</lparam></gate>
<gate>
<ID>258</ID>
<type>DE_TO</type>
<position>309.5,-194.5</position>
<input>
<ID>IN_0</ID>976 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_ACC_OUT</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_LABEL</type>
<position>211,8</position>
<gparam>LABEL_TEXT PROCESSADOR BIP IMT - MAUA 2022</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>1048</ID>
<type>DE_TO</type>
<position>253,-98</position>
<input>
<ID>IN_0</ID>283 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_ACC_IN</lparam></gate>
<gate>
<ID>1049</ID>
<type>DE_TO</type>
<position>253.5,-110</position>
<input>
<ID>IN_0</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_ACC_IN</lparam></gate>
<gate>
<ID>1050</ID>
<type>DE_TO</type>
<position>254,-122.5</position>
<input>
<ID>IN_0</ID>295 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_ACC_IN</lparam></gate>
<gate>
<ID>1051</ID>
<type>DE_TO</type>
<position>255.5,-135.5</position>
<input>
<ID>IN_0</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_ACC_IN</lparam></gate>
<gate>
<ID>1052</ID>
<type>DE_TO</type>
<position>254.5,-149</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_ACC_IN</lparam></gate>
<gate>
<ID>1053</ID>
<type>DE_TO</type>
<position>254.5,-162</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_ACC_IN</lparam></gate>
<gate>
<ID>1054</ID>
<type>DE_TO</type>
<position>254,-175</position>
<input>
<ID>IN_0</ID>319 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_ACC_IN</lparam></gate>
<gate>
<ID>1055</ID>
<type>DE_TO</type>
<position>254.5,-189</position>
<input>
<ID>IN_0</ID>325 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_ACC_IN</lparam></gate>
<gate>
<ID>1056</ID>
<type>DE_TO</type>
<position>255,-203</position>
<input>
<ID>IN_0</ID>331 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_ACC_IN</lparam></gate>
<gate>
<ID>1057</ID>
<type>DE_TO</type>
<position>254,-216</position>
<input>
<ID>IN_0</ID>337 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_ACC_IN</lparam></gate>
<gate>
<ID>1058</ID>
<type>DE_TO</type>
<position>254.5,-229</position>
<input>
<ID>IN_0</ID>343 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_ACC_IN</lparam></gate>
<gate>
<ID>1059</ID>
<type>DE_TO</type>
<position>253.5,-242.5</position>
<input>
<ID>IN_0</ID>349 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_ACC_IN</lparam></gate>
<gate>
<ID>291</ID>
<type>DA_FROM</type>
<position>270.5,-54.5</position>
<input>
<ID>IN_0</ID>210 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RESET</lparam></gate>
<gate>
<ID>304</ID>
<type>DE_TO</type>
<position>309.5,-208.5</position>
<input>
<ID>IN_0</ID>978 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_ACC_OUT</lparam></gate>
<gate>
<ID>305</ID>
<type>DE_TO</type>
<position>309,-221.5</position>
<input>
<ID>IN_0</ID>980 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_ACC_OUT</lparam></gate>
<gate>
<ID>306</ID>
<type>DE_TO</type>
<position>309,-234.5</position>
<input>
<ID>IN_0</ID>982 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_ACC_OUT</lparam></gate>
<gate>
<ID>307</ID>
<type>DE_TO</type>
<position>309.5,-248.5</position>
<input>
<ID>IN_0</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_ACC_OUT</lparam></gate>
<gate>
<ID>317</ID>
<type>DA_FROM</type>
<position>207.5,-45.5</position>
<input>
<ID>IN_0</ID>255 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>319</ID>
<type>DA_FROM</type>
<position>207.5,-42.5</position>
<input>
<ID>IN_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>321</ID>
<type>DA_FROM</type>
<position>222.5,-54.5</position>
<input>
<ID>IN_0</ID>257 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_RAM</lparam></gate>
<gate>
<ID>323</ID>
<type>DA_FROM</type>
<position>211.5,-52.5</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_ES</lparam></gate>
<gate>
<ID>325</ID>
<type>DA_FROM</type>
<position>203,-50.5</position>
<input>
<ID>IN_0</ID>259 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_ULA</lparam></gate>
<gate>
<ID>326</ID>
<type>AE_MUX_4x1</type>
<position>186,-64.5</position>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>263 </input>
<input>
<ID>IN_2</ID>264 </input>
<output>
<ID>OUT</ID>265 </output>
<input>
<ID>SEL_0</ID>261 </input>
<input>
<ID>SEL_1</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>327</ID>
<type>DA_FROM</type>
<position>165,-58.5</position>
<input>
<ID>IN_0</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>328</ID>
<type>DA_FROM</type>
<position>165,-55.5</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>329</ID>
<type>DA_FROM</type>
<position>179.5,-67.5</position>
<input>
<ID>IN_0</ID>262 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_RAM</lparam></gate>
<gate>
<ID>330</ID>
<type>DA_FROM</type>
<position>168.5,-65.5</position>
<input>
<ID>IN_0</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_ES</lparam></gate>
<gate>
<ID>331</ID>
<type>DA_FROM</type>
<position>160,-63.5</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_ULA</lparam></gate>
<gate>
<ID>332</ID>
<type>AE_MUX_4x1</type>
<position>229.5,-77.5</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>269 </input>
<input>
<ID>IN_2</ID>270 </input>
<output>
<ID>OUT</ID>271 </output>
<input>
<ID>SEL_0</ID>267 </input>
<input>
<ID>SEL_1</ID>266 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>333</ID>
<type>DA_FROM</type>
<position>208.5,-71.5</position>
<input>
<ID>IN_0</ID>266 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>1112</ID>
<type>AA_LABEL</type>
<position>228.5,-23</position>
<gparam>LABEL_TEXT Acumulador</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>334</ID>
<type>DA_FROM</type>
<position>208.5,-68.5</position>
<input>
<ID>IN_0</ID>267 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>335</ID>
<type>DA_FROM</type>
<position>223,-80.5</position>
<input>
<ID>IN_0</ID>268 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_RAM</lparam></gate>
<gate>
<ID>336</ID>
<type>DA_FROM</type>
<position>212,-78.5</position>
<input>
<ID>IN_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_ES</lparam></gate>
<gate>
<ID>337</ID>
<type>DA_FROM</type>
<position>203.5,-76.5</position>
<input>
<ID>IN_0</ID>270 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_ULA</lparam></gate>
<gate>
<ID>338</ID>
<type>AE_MUX_4x1</type>
<position>185.5,-90.5</position>
<input>
<ID>IN_0</ID>274 </input>
<input>
<ID>IN_1</ID>275 </input>
<input>
<ID>IN_2</ID>276 </input>
<output>
<ID>OUT</ID>277 </output>
<input>
<ID>SEL_0</ID>273 </input>
<input>
<ID>SEL_1</ID>272 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>339</ID>
<type>DA_FROM</type>
<position>164.5,-84.5</position>
<input>
<ID>IN_0</ID>272 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>340</ID>
<type>DA_FROM</type>
<position>164.5,-81.5</position>
<input>
<ID>IN_0</ID>273 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>341</ID>
<type>DA_FROM</type>
<position>179,-93.5</position>
<input>
<ID>IN_0</ID>274 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_RAM</lparam></gate>
<gate>
<ID>342</ID>
<type>DA_FROM</type>
<position>168,-91.5</position>
<input>
<ID>IN_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_ES</lparam></gate>
<gate>
<ID>343</ID>
<type>DA_FROM</type>
<position>159.5,-89.5</position>
<input>
<ID>IN_0</ID>276 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_ULA</lparam></gate>
<gate>
<ID>344</ID>
<type>AE_MUX_4x1</type>
<position>230.5,-103.5</position>
<input>
<ID>IN_0</ID>280 </input>
<input>
<ID>IN_1</ID>281 </input>
<input>
<ID>IN_2</ID>282 </input>
<output>
<ID>OUT</ID>283 </output>
<input>
<ID>SEL_0</ID>279 </input>
<input>
<ID>SEL_1</ID>278 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>345</ID>
<type>DA_FROM</type>
<position>209.5,-97.5</position>
<input>
<ID>IN_0</ID>278 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>346</ID>
<type>DA_FROM</type>
<position>209.5,-94.5</position>
<input>
<ID>IN_0</ID>279 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>347</ID>
<type>DA_FROM</type>
<position>224,-106.5</position>
<input>
<ID>IN_0</ID>280 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_RAM</lparam></gate>
<gate>
<ID>348</ID>
<type>DA_FROM</type>
<position>213,-104.5</position>
<input>
<ID>IN_0</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_ES</lparam></gate>
<gate>
<ID>349</ID>
<type>DA_FROM</type>
<position>204.5,-102.5</position>
<input>
<ID>IN_0</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_ULA</lparam></gate>
<gate>
<ID>350</ID>
<type>AE_MUX_4x1</type>
<position>186,-115.5</position>
<input>
<ID>IN_0</ID>286 </input>
<input>
<ID>IN_1</ID>287 </input>
<input>
<ID>IN_2</ID>288 </input>
<output>
<ID>OUT</ID>289 </output>
<input>
<ID>SEL_0</ID>285 </input>
<input>
<ID>SEL_1</ID>284 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>351</ID>
<type>DA_FROM</type>
<position>163.5,-109.5</position>
<input>
<ID>IN_0</ID>284 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>352</ID>
<type>DA_FROM</type>
<position>163.5,-106.5</position>
<input>
<ID>IN_0</ID>285 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>353</ID>
<type>DA_FROM</type>
<position>178,-118.5</position>
<input>
<ID>IN_0</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_RAM</lparam></gate>
<gate>
<ID>1132</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>412.5,-67.5</position>
<input>
<ID>IN_0</ID>911 </input>
<input>
<ID>IN_1</ID>912 </input>
<input>
<ID>IN_2</ID>913 </input>
<input>
<ID>IN_3</ID>914 </input>
<input>
<ID>IN_4</ID>910 </input>
<input>
<ID>IN_5</ID>909 </input>
<input>
<ID>IN_6</ID>908 </input>
<input>
<ID>IN_7</ID>907 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 49</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>354</ID>
<type>DA_FROM</type>
<position>167,-116.5</position>
<input>
<ID>IN_0</ID>287 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_ES</lparam></gate>
<gate>
<ID>1133</ID>
<type>DA_FROM</type>
<position>406,-59</position>
<input>
<ID>IN_0</ID>907 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D7_ACC_IN</lparam></gate>
<gate>
<ID>355</ID>
<type>DA_FROM</type>
<position>158.5,-114.5</position>
<input>
<ID>IN_0</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_ULA</lparam></gate>
<gate>
<ID>1134</ID>
<type>DA_FROM</type>
<position>407.5,-56</position>
<input>
<ID>IN_0</ID>908 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D6_ACC_IN</lparam></gate>
<gate>
<ID>356</ID>
<type>AE_MUX_4x1</type>
<position>230.5,-128.5</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>293 </input>
<input>
<ID>IN_2</ID>294 </input>
<output>
<ID>OUT</ID>295 </output>
<input>
<ID>SEL_0</ID>291 </input>
<input>
<ID>SEL_1</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1135</ID>
<type>DA_FROM</type>
<position>406,-53</position>
<input>
<ID>IN_0</ID>909 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D5_ACC_IN</lparam></gate>
<gate>
<ID>357</ID>
<type>DA_FROM</type>
<position>209.5,-122.5</position>
<input>
<ID>IN_0</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>1136</ID>
<type>DA_FROM</type>
<position>406,-50</position>
<input>
<ID>IN_0</ID>910 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D4_ACC_IN</lparam></gate>
<gate>
<ID>358</ID>
<type>DA_FROM</type>
<position>209.5,-119.5</position>
<input>
<ID>IN_0</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>1137</ID>
<type>DA_FROM</type>
<position>406,-84</position>
<input>
<ID>IN_0</ID>914 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D3_ACC_IN</lparam></gate>
<gate>
<ID>359</ID>
<type>DA_FROM</type>
<position>224,-131.5</position>
<input>
<ID>IN_0</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_RAM</lparam></gate>
<gate>
<ID>1138</ID>
<type>DA_FROM</type>
<position>406,-81</position>
<input>
<ID>IN_0</ID>913 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D2_ACC_IN</lparam></gate>
<gate>
<ID>360</ID>
<type>DA_FROM</type>
<position>213,-129.5</position>
<input>
<ID>IN_0</ID>293 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_ES</lparam></gate>
<gate>
<ID>1139</ID>
<type>DA_FROM</type>
<position>406,-78</position>
<input>
<ID>IN_0</ID>912 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D1_ACC_IN</lparam></gate>
<gate>
<ID>361</ID>
<type>DA_FROM</type>
<position>204.5,-127.5</position>
<input>
<ID>IN_0</ID>294 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_ULA</lparam></gate>
<gate>
<ID>1140</ID>
<type>DA_FROM</type>
<position>406,-75</position>
<input>
<ID>IN_0</ID>911 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D0_ACC_IN</lparam></gate>
<gate>
<ID>362</ID>
<type>AE_MUX_4x1</type>
<position>187,-141.5</position>
<input>
<ID>IN_0</ID>298 </input>
<input>
<ID>IN_1</ID>299 </input>
<input>
<ID>IN_2</ID>300 </input>
<output>
<ID>OUT</ID>301 </output>
<input>
<ID>SEL_0</ID>297 </input>
<input>
<ID>SEL_1</ID>296 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1141</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>389,-67</position>
<input>
<ID>IN_0</ID>919 </input>
<input>
<ID>IN_1</ID>920 </input>
<input>
<ID>IN_2</ID>921 </input>
<input>
<ID>IN_3</ID>922 </input>
<input>
<ID>IN_4</ID>918 </input>
<input>
<ID>IN_5</ID>917 </input>
<input>
<ID>IN_6</ID>916 </input>
<input>
<ID>IN_7</ID>915 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 218</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>363</ID>
<type>DA_FROM</type>
<position>166,-135.5</position>
<input>
<ID>IN_0</ID>296 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>1142</ID>
<type>DA_FROM</type>
<position>382.5,-58.5</position>
<input>
<ID>IN_0</ID>915 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D15_ACC_IN</lparam></gate>
<gate>
<ID>364</ID>
<type>DA_FROM</type>
<position>166,-132.5</position>
<input>
<ID>IN_0</ID>297 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>1143</ID>
<type>DA_FROM</type>
<position>382.5,-55.5</position>
<input>
<ID>IN_0</ID>916 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D14_ACC_IN</lparam></gate>
<gate>
<ID>365</ID>
<type>DA_FROM</type>
<position>180.5,-144.5</position>
<input>
<ID>IN_0</ID>298 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_RAM</lparam></gate>
<gate>
<ID>1144</ID>
<type>DA_FROM</type>
<position>382.5,-52.5</position>
<input>
<ID>IN_0</ID>917 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D13_ACC_IN</lparam></gate>
<gate>
<ID>366</ID>
<type>DA_FROM</type>
<position>169.5,-142.5</position>
<input>
<ID>IN_0</ID>299 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_ES</lparam></gate>
<gate>
<ID>1145</ID>
<type>DA_FROM</type>
<position>382.5,-49.5</position>
<input>
<ID>IN_0</ID>918 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D12_ACC_IN</lparam></gate>
<gate>
<ID>367</ID>
<type>DA_FROM</type>
<position>161,-140.5</position>
<input>
<ID>IN_0</ID>300 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_ULA</lparam></gate>
<gate>
<ID>1146</ID>
<type>DA_FROM</type>
<position>382.5,-83.5</position>
<input>
<ID>IN_0</ID>922 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D11_ACC_IN</lparam></gate>
<gate>
<ID>368</ID>
<type>AE_MUX_4x1</type>
<position>231.5,-154.5</position>
<input>
<ID>IN_0</ID>304 </input>
<input>
<ID>IN_1</ID>305 </input>
<input>
<ID>IN_2</ID>306 </input>
<output>
<ID>OUT</ID>307 </output>
<input>
<ID>SEL_0</ID>303 </input>
<input>
<ID>SEL_1</ID>302 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1147</ID>
<type>DA_FROM</type>
<position>382.5,-80.5</position>
<input>
<ID>IN_0</ID>921 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D10_ACC_IN</lparam></gate>
<gate>
<ID>369</ID>
<type>DA_FROM</type>
<position>210.5,-148.5</position>
<input>
<ID>IN_0</ID>302 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>1148</ID>
<type>DA_FROM</type>
<position>382.5,-77.5</position>
<input>
<ID>IN_0</ID>920 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D9_ACC_IN</lparam></gate>
<gate>
<ID>370</ID>
<type>DA_FROM</type>
<position>210.5,-145.5</position>
<input>
<ID>IN_0</ID>303 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>1149</ID>
<type>DA_FROM</type>
<position>382.5,-74.5</position>
<input>
<ID>IN_0</ID>919 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D8_ACC_IN</lparam></gate>
<gate>
<ID>371</ID>
<type>DA_FROM</type>
<position>225,-157.5</position>
<input>
<ID>IN_0</ID>304 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_RAM</lparam></gate>
<gate>
<ID>1150</ID>
<type>AA_LABEL</type>
<position>397,-38.5</position>
<gparam>LABEL_TEXT Acumulador IN</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>372</ID>
<type>DA_FROM</type>
<position>214,-155.5</position>
<input>
<ID>IN_0</ID>305 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_ES</lparam></gate>
<gate>
<ID>373</ID>
<type>DA_FROM</type>
<position>205.5,-153.5</position>
<input>
<ID>IN_0</ID>306 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_ULA</lparam></gate>
<gate>
<ID>374</ID>
<type>AE_MUX_4x1</type>
<position>187.5,-167.5</position>
<input>
<ID>IN_0</ID>310 </input>
<input>
<ID>IN_1</ID>311 </input>
<input>
<ID>IN_2</ID>312 </input>
<output>
<ID>OUT</ID>313 </output>
<input>
<ID>SEL_0</ID>309 </input>
<input>
<ID>SEL_1</ID>308 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>375</ID>
<type>DA_FROM</type>
<position>166.5,-161.5</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>376</ID>
<type>DA_FROM</type>
<position>166.5,-158.5</position>
<input>
<ID>IN_0</ID>309 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>377</ID>
<type>DA_FROM</type>
<position>181,-170.5</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_RAM</lparam></gate>
<gate>
<ID>378</ID>
<type>DA_FROM</type>
<position>170,-168.5</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_ES</lparam></gate>
<gate>
<ID>379</ID>
<type>DA_FROM</type>
<position>161.5,-166.5</position>
<input>
<ID>IN_0</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_ULA</lparam></gate>
<gate>
<ID>380</ID>
<type>AE_MUX_4x1</type>
<position>233.5,-180.5</position>
<input>
<ID>IN_0</ID>316 </input>
<input>
<ID>IN_1</ID>317 </input>
<input>
<ID>IN_2</ID>318 </input>
<output>
<ID>OUT</ID>319 </output>
<input>
<ID>SEL_0</ID>315 </input>
<input>
<ID>SEL_1</ID>314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>381</ID>
<type>DA_FROM</type>
<position>212,-174.5</position>
<input>
<ID>IN_0</ID>314 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>382</ID>
<type>DA_FROM</type>
<position>212,-171.5</position>
<input>
<ID>IN_0</ID>315 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>383</ID>
<type>DA_FROM</type>
<position>226.5,-183.5</position>
<input>
<ID>IN_0</ID>316 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_RAM</lparam></gate>
<gate>
<ID>384</ID>
<type>DA_FROM</type>
<position>215.5,-181.5</position>
<input>
<ID>IN_0</ID>317 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_ES</lparam></gate>
<gate>
<ID>385</ID>
<type>DA_FROM</type>
<position>207,-179.5</position>
<input>
<ID>IN_0</ID>318 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_ULA</lparam></gate>
<gate>
<ID>386</ID>
<type>AE_MUX_4x1</type>
<position>188.5,-194.5</position>
<input>
<ID>IN_0</ID>322 </input>
<input>
<ID>IN_1</ID>323 </input>
<input>
<ID>IN_2</ID>324 </input>
<output>
<ID>OUT</ID>325 </output>
<input>
<ID>SEL_0</ID>321 </input>
<input>
<ID>SEL_1</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>387</ID>
<type>DA_FROM</type>
<position>167.5,-188.5</position>
<input>
<ID>IN_0</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<gate>
<ID>388</ID>
<type>DA_FROM</type>
<position>167.5,-185.5</position>
<input>
<ID>IN_0</ID>321 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<wire>
<ID>965</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-128,294.5,-128</points>
<connection>
<GID>1200</GID>
<name>clock</name></connection>
<connection>
<GID>1199</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>966</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,-128.5,303.5,-126</points>
<intersection>-128.5 1</intersection>
<intersection>-126 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-128.5,307,-128.5</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300.5,-126,303.5,-126</points>
<connection>
<GID>1200</GID>
<name>OUT_0</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>967</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290.5,-142,295,-142</points>
<connection>
<GID>1202</GID>
<name>clock</name></connection>
<connection>
<GID>1201</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>968</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,-141.5,304,-140</points>
<intersection>-141.5 1</intersection>
<intersection>-140 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-141.5,307,-141.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>304 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,-140,304,-140</points>
<connection>
<GID>1202</GID>
<name>OUT_0</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>969</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290.5,-155,295,-155</points>
<connection>
<GID>1204</GID>
<name>clock</name></connection>
<connection>
<GID>1203</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>970</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,-154.5,304,-153</points>
<intersection>-154.5 1</intersection>
<intersection>-153 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-154.5,307.5,-154.5</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>304 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,-153,304,-153</points>
<connection>
<GID>1204</GID>
<name>OUT_0</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>971</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290.5,-167.5,295,-167.5</points>
<connection>
<GID>1206</GID>
<name>clock</name></connection>
<connection>
<GID>1205</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>972</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,-167.5,304,-165.5</points>
<intersection>-167.5 1</intersection>
<intersection>-165.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-167.5,307.5,-167.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>304 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,-165.5,304,-165.5</points>
<connection>
<GID>1206</GID>
<name>OUT_0</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>973</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-181.5,294.5,-181.5</points>
<connection>
<GID>1208</GID>
<name>clock</name></connection>
<connection>
<GID>1207</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>974</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,-180.5,303.5,-179.5</points>
<intersection>-180.5 1</intersection>
<intersection>-179.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-180.5,307,-180.5</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300.5,-179.5,303.5,-179.5</points>
<connection>
<GID>1208</GID>
<name>OUT_0</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>975</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290.5,-195.5,294.5,-195.5</points>
<connection>
<GID>1210</GID>
<name>clock</name></connection>
<connection>
<GID>1209</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>976</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,-194.5,304.5,-193.5</points>
<intersection>-194.5 1</intersection>
<intersection>-193.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,-194.5,307.5,-194.5</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300.5,-193.5,304.5,-193.5</points>
<connection>
<GID>1210</GID>
<name>OUT_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>977</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289.5,-208.5,294,-208.5</points>
<connection>
<GID>1212</GID>
<name>clock</name></connection>
<connection>
<GID>1211</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>978</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,-208.5,303.5,-206.5</points>
<intersection>-208.5 1</intersection>
<intersection>-206.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-208.5,307.5,-208.5</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300,-206.5,303.5,-206.5</points>
<connection>
<GID>1212</GID>
<name>OUT_0</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>979</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-221,294,-221</points>
<connection>
<GID>1214</GID>
<name>clock</name></connection>
<connection>
<GID>1213</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>980</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,-221.5,303.5,-219</points>
<intersection>-221.5 1</intersection>
<intersection>-219 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-221.5,307,-221.5</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300,-219,303.5,-219</points>
<connection>
<GID>1214</GID>
<name>OUT_0</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>981</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289.5,-235,294,-235</points>
<connection>
<GID>1216</GID>
<name>clock</name></connection>
<connection>
<GID>1215</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>272.5,-51.5,278.5,-51.5</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>278.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>278.5,-251,278.5,-51.5</points>
<intersection>-251 117</intersection>
<intersection>-237 115</intersection>
<intersection>-223 113</intersection>
<intersection>-210.5 111</intersection>
<intersection>-197.5 109</intersection>
<intersection>-183.5 107</intersection>
<intersection>-169.5 105</intersection>
<intersection>-157 103</intersection>
<intersection>-144 101</intersection>
<intersection>-130 99</intersection>
<intersection>-117.5 97</intersection>
<intersection>-105.5 95</intersection>
<intersection>-93.5 93</intersection>
<intersection>-80 91</intersection>
<intersection>-67.5 89</intersection>
<intersection>-55.5 87</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>87</ID>
<points>278.5,-55.5,296,-55.5</points>
<connection>
<GID>1186</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>89</ID>
<points>278.5,-67.5,296.5,-67.5</points>
<connection>
<GID>1190</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>91</ID>
<points>278.5,-80,294.5,-80</points>
<connection>
<GID>1192</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>93</ID>
<points>278.5,-93.5,294.5,-93.5</points>
<connection>
<GID>1194</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>95</ID>
<points>278.5,-105.5,295,-105.5</points>
<connection>
<GID>1196</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>97</ID>
<points>278.5,-117.5,294.5,-117.5</points>
<connection>
<GID>1198</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>99</ID>
<points>278.5,-130,294.5,-130</points>
<connection>
<GID>1200</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>101</ID>
<points>278.5,-144,295,-144</points>
<connection>
<GID>1202</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>103</ID>
<points>278.5,-157,295,-157</points>
<connection>
<GID>1204</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>105</ID>
<points>278.5,-169.5,295,-169.5</points>
<connection>
<GID>1206</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>107</ID>
<points>278.5,-183.5,294.5,-183.5</points>
<connection>
<GID>1208</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>109</ID>
<points>278.5,-197.5,294.5,-197.5</points>
<connection>
<GID>1210</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>111</ID>
<points>278.5,-210.5,294,-210.5</points>
<connection>
<GID>1212</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>113</ID>
<points>278.5,-223,294,-223</points>
<connection>
<GID>1214</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>115</ID>
<points>278.5,-237,294,-237</points>
<connection>
<GID>1216</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment>
<hsegment>
<ID>117</ID>
<points>278.5,-251,294.5,-251</points>
<connection>
<GID>1218</GID>
<name>clock_enable</name></connection>
<intersection>278.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>982</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,-234.5,303.5,-233</points>
<intersection>-234.5 1</intersection>
<intersection>-233 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-234.5,307,-234.5</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300,-233,303.5,-233</points>
<connection>
<GID>1216</GID>
<name>OUT_0</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>272.5,-54.5,275.5,-54.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>275.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>275.5,-254,275.5,-54.5</points>
<intersection>-254 149</intersection>
<intersection>-240 147</intersection>
<intersection>-226.5 144</intersection>
<intersection>-213 141</intersection>
<intersection>-201 138</intersection>
<intersection>-187 135</intersection>
<intersection>-172.5 132</intersection>
<intersection>-160 129</intersection>
<intersection>-147 126</intersection>
<intersection>-133.5 122</intersection>
<intersection>-121 121</intersection>
<intersection>-109 115</intersection>
<intersection>-97 112</intersection>
<intersection>-83 109</intersection>
<intersection>-71 105</intersection>
<intersection>-58.5 102</intersection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>102</ID>
<points>275.5,-58.5,299,-58.5</points>
<intersection>275.5 2</intersection>
<intersection>299 107</intersection></hsegment>
<hsegment>
<ID>105</ID>
<points>275.5,-71,299.5,-71</points>
<intersection>275.5 2</intersection>
<intersection>299.5 106</intersection></hsegment>
<vsegment>
<ID>106</ID>
<points>299.5,-71,299.5,-69.5</points>
<connection>
<GID>1190</GID>
<name>clear</name></connection>
<intersection>-71 105</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>299,-58.5,299,-57.5</points>
<connection>
<GID>1186</GID>
<name>clear</name></connection>
<intersection>-58.5 102</intersection></vsegment>
<hsegment>
<ID>109</ID>
<points>275.5,-83,297.5,-83</points>
<intersection>275.5 2</intersection>
<intersection>297.5 110</intersection></hsegment>
<vsegment>
<ID>110</ID>
<points>297.5,-83,297.5,-82</points>
<connection>
<GID>1192</GID>
<name>clear</name></connection>
<intersection>-83 109</intersection></vsegment>
<hsegment>
<ID>112</ID>
<points>275.5,-97,297.5,-97</points>
<intersection>275.5 2</intersection>
<intersection>297.5 113</intersection></hsegment>
<vsegment>
<ID>113</ID>
<points>297.5,-97,297.5,-95.5</points>
<connection>
<GID>1194</GID>
<name>clear</name></connection>
<intersection>-97 112</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>275.5,-109,298,-109</points>
<intersection>275.5 2</intersection>
<intersection>298 116</intersection></hsegment>
<vsegment>
<ID>116</ID>
<points>298,-109,298,-107.5</points>
<connection>
<GID>1196</GID>
<name>clear</name></connection>
<intersection>-109 115</intersection></vsegment>
<hsegment>
<ID>121</ID>
<points>275.5,-121,297.5,-121</points>
<intersection>275.5 2</intersection>
<intersection>297.5 124</intersection></hsegment>
<hsegment>
<ID>122</ID>
<points>275.5,-133.5,297.5,-133.5</points>
<intersection>275.5 2</intersection>
<intersection>297.5 123</intersection></hsegment>
<vsegment>
<ID>123</ID>
<points>297.5,-133.5,297.5,-132</points>
<connection>
<GID>1200</GID>
<name>clear</name></connection>
<intersection>-133.5 122</intersection></vsegment>
<vsegment>
<ID>124</ID>
<points>297.5,-121,297.5,-119.5</points>
<connection>
<GID>1198</GID>
<name>clear</name></connection>
<intersection>-121 121</intersection></vsegment>
<hsegment>
<ID>126</ID>
<points>275.5,-147,298,-147</points>
<intersection>275.5 2</intersection>
<intersection>298 127</intersection></hsegment>
<vsegment>
<ID>127</ID>
<points>298,-147,298,-146</points>
<connection>
<GID>1202</GID>
<name>clear</name></connection>
<intersection>-147 126</intersection></vsegment>
<hsegment>
<ID>129</ID>
<points>275.5,-160,298,-160</points>
<intersection>275.5 2</intersection>
<intersection>298 130</intersection></hsegment>
<vsegment>
<ID>130</ID>
<points>298,-160,298,-159</points>
<connection>
<GID>1204</GID>
<name>clear</name></connection>
<intersection>-160 129</intersection></vsegment>
<hsegment>
<ID>132</ID>
<points>275.5,-172.5,298,-172.5</points>
<intersection>275.5 2</intersection>
<intersection>298 133</intersection></hsegment>
<vsegment>
<ID>133</ID>
<points>298,-172.5,298,-171.5</points>
<connection>
<GID>1206</GID>
<name>clear</name></connection>
<intersection>-172.5 132</intersection></vsegment>
<hsegment>
<ID>135</ID>
<points>275.5,-187,297.5,-187</points>
<intersection>275.5 2</intersection>
<intersection>297.5 136</intersection></hsegment>
<vsegment>
<ID>136</ID>
<points>297.5,-187,297.5,-185.5</points>
<connection>
<GID>1208</GID>
<name>clear</name></connection>
<intersection>-187 135</intersection></vsegment>
<hsegment>
<ID>138</ID>
<points>275.5,-201,297.5,-201</points>
<intersection>275.5 2</intersection>
<intersection>297.5 139</intersection></hsegment>
<vsegment>
<ID>139</ID>
<points>297.5,-201,297.5,-199.5</points>
<connection>
<GID>1210</GID>
<name>clear</name></connection>
<intersection>-201 138</intersection></vsegment>
<hsegment>
<ID>141</ID>
<points>275.5,-213,297,-213</points>
<intersection>275.5 2</intersection>
<intersection>297 142</intersection></hsegment>
<vsegment>
<ID>142</ID>
<points>297,-213,297,-212.5</points>
<connection>
<GID>1212</GID>
<name>clear</name></connection>
<intersection>-213 141</intersection></vsegment>
<hsegment>
<ID>144</ID>
<points>275.5,-226.5,297,-226.5</points>
<intersection>275.5 2</intersection>
<intersection>297 145</intersection></hsegment>
<vsegment>
<ID>145</ID>
<points>297,-226.5,297,-225</points>
<connection>
<GID>1214</GID>
<name>clear</name></connection>
<intersection>-226.5 144</intersection></vsegment>
<hsegment>
<ID>147</ID>
<points>275.5,-240,297,-240</points>
<intersection>275.5 2</intersection>
<intersection>297 150</intersection></hsegment>
<hsegment>
<ID>149</ID>
<points>275.5,-254,297.5,-254</points>
<intersection>275.5 2</intersection>
<intersection>297.5 151</intersection></hsegment>
<vsegment>
<ID>150</ID>
<points>297,-240,297,-239</points>
<connection>
<GID>1216</GID>
<name>clear</name></connection>
<intersection>-240 147</intersection></vsegment>
<vsegment>
<ID>151</ID>
<points>297.5,-254,297.5,-253</points>
<connection>
<GID>1218</GID>
<name>clear</name></connection>
<intersection>-254 149</intersection></vsegment></shape></wire>
<wire>
<ID>983</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-249,294.5,-249</points>
<connection>
<GID>1218</GID>
<name>clock</name></connection>
<connection>
<GID>1217</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>984</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,-248.5,304,-247</points>
<intersection>-248.5 1</intersection>
<intersection>-247 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-248.5,307.5,-248.5</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>304 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300.5,-247,304,-247</points>
<connection>
<GID>1218</GID>
<name>OUT_0</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-46.5,229,-45.5</points>
<connection>
<GID>246</GID>
<name>SEL_1</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>209.5,-45.5,229,-45.5</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-46.5,230,-42.5</points>
<connection>
<GID>246</GID>
<name>SEL_0</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>209.5,-42.5,230,-42.5</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>224.5,-54.5,226,-54.5</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<connection>
<GID>321</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213.5,-52.5,226,-52.5</points>
<connection>
<GID>246</GID>
<name>IN_1</name></connection>
<connection>
<GID>323</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>205,-50.5,226,-50.5</points>
<connection>
<GID>246</GID>
<name>IN_2</name></connection>
<connection>
<GID>325</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,-59.5,186,-58.5</points>
<connection>
<GID>326</GID>
<name>SEL_1</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,-58.5,186,-58.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>186 0</intersection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187,-59.5,187,-55.5</points>
<connection>
<GID>326</GID>
<name>SEL_0</name></connection>
<intersection>-55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,-55.5,187,-55.5</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>181.5,-67.5,183,-67.5</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<connection>
<GID>329</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170.5,-65.5,183,-65.5</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<connection>
<GID>330</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-63.5,183,-63.5</points>
<connection>
<GID>326</GID>
<name>IN_2</name></connection>
<connection>
<GID>331</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189,-64.5,239.5,-64.5</points>
<connection>
<GID>326</GID>
<name>OUT</name></connection>
<intersection>239.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>239.5,-64.5,239.5,-59</points>
<connection>
<GID>1025</GID>
<name>IN_0</name></connection>
<intersection>-64.5 1</intersection>
<intersection>-63.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>239.5,-63.5,296.5,-63.5</points>
<connection>
<GID>1190</GID>
<name>IN_0</name></connection>
<intersection>239.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,-72.5,229.5,-71.5</points>
<connection>
<GID>332</GID>
<name>SEL_1</name></connection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>210.5,-71.5,229.5,-71.5</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>229.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-72.5,230.5,-68.5</points>
<connection>
<GID>332</GID>
<name>SEL_0</name></connection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>210.5,-68.5,230.5,-68.5</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<intersection>230.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-80.5,226.5,-80.5</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<connection>
<GID>335</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>214,-78.5,226.5,-78.5</points>
<connection>
<GID>332</GID>
<name>IN_1</name></connection>
<connection>
<GID>336</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>205.5,-76.5,226.5,-76.5</points>
<connection>
<GID>332</GID>
<name>IN_2</name></connection>
<connection>
<GID>337</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>232.5,-77.5,249.5,-77.5</points>
<connection>
<GID>332</GID>
<name>OUT</name></connection>
<intersection>249.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>249.5,-77.5,249.5,-71</points>
<connection>
<GID>1026</GID>
<name>IN_0</name></connection>
<intersection>-77.5 1</intersection>
<intersection>-76 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>249.5,-76,294.5,-76</points>
<connection>
<GID>1192</GID>
<name>IN_0</name></connection>
<intersection>249.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-85.5,185.5,-84.5</points>
<connection>
<GID>338</GID>
<name>SEL_1</name></connection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,-84.5,185.5,-84.5</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,-85.5,186.5,-81.5</points>
<connection>
<GID>338</GID>
<name>SEL_0</name></connection>
<intersection>-81.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,-81.5,186.5,-81.5</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>181,-93.5,182.5,-93.5</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<connection>
<GID>341</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-91.5,182.5,-91.5</points>
<connection>
<GID>338</GID>
<name>IN_1</name></connection>
<connection>
<GID>342</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,-89.5,182.5,-89.5</points>
<connection>
<GID>338</GID>
<name>IN_2</name></connection>
<connection>
<GID>343</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>188.5,-90.5,249,-90.5</points>
<connection>
<GID>338</GID>
<name>OUT</name></connection>
<intersection>249 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>249,-90.5,249,-84</points>
<connection>
<GID>1027</GID>
<name>IN_0</name></connection>
<intersection>-90.5 1</intersection>
<intersection>-89.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>249,-89.5,294.5,-89.5</points>
<connection>
<GID>1194</GID>
<name>IN_0</name></connection>
<intersection>249 2</intersection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-98.5,230.5,-97.5</points>
<connection>
<GID>344</GID>
<name>SEL_1</name></connection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211.5,-97.5,230.5,-97.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>230.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-98.5,231.5,-94.5</points>
<connection>
<GID>344</GID>
<name>SEL_0</name></connection>
<intersection>-94.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211.5,-94.5,231.5,-94.5</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>231.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>226,-106.5,227.5,-106.5</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<connection>
<GID>347</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215,-104.5,227.5,-104.5</points>
<connection>
<GID>344</GID>
<name>IN_1</name></connection>
<connection>
<GID>348</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>206.5,-102.5,227.5,-102.5</points>
<connection>
<GID>344</GID>
<name>IN_2</name></connection>
<connection>
<GID>349</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>233.5,-103.5,251,-103.5</points>
<connection>
<GID>344</GID>
<name>OUT</name></connection>
<intersection>251 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>251,-103.5,251,-98</points>
<connection>
<GID>1048</GID>
<name>IN_0</name></connection>
<intersection>-103.5 1</intersection>
<intersection>-101.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>251,-101.5,295,-101.5</points>
<connection>
<GID>1196</GID>
<name>IN_0</name></connection>
<intersection>251 2</intersection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,-110.5,186,-109.5</points>
<connection>
<GID>350</GID>
<name>SEL_1</name></connection>
<intersection>-109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165.5,-109.5,186,-109.5</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>186 0</intersection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187,-110.5,187,-106.5</points>
<connection>
<GID>350</GID>
<name>SEL_0</name></connection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165.5,-106.5,187,-106.5</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>180,-118.5,183,-118.5</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<connection>
<GID>353</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-116.5,183,-116.5</points>
<connection>
<GID>350</GID>
<name>IN_1</name></connection>
<connection>
<GID>354</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>160.5,-114.5,183,-114.5</points>
<connection>
<GID>350</GID>
<name>IN_2</name></connection>
<connection>
<GID>355</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189,-115.5,251.5,-115.5</points>
<connection>
<GID>350</GID>
<name>OUT</name></connection>
<intersection>251.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>251.5,-115.5,251.5,-110</points>
<connection>
<GID>1049</GID>
<name>IN_0</name></connection>
<intersection>-115.5 1</intersection>
<intersection>-113.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>251.5,-113.5,294.5,-113.5</points>
<connection>
<GID>1198</GID>
<name>IN_0</name></connection>
<intersection>251.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-123.5,230.5,-122.5</points>
<connection>
<GID>356</GID>
<name>SEL_1</name></connection>
<intersection>-122.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211.5,-122.5,230.5,-122.5</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<intersection>230.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-123.5,231.5,-119.5</points>
<connection>
<GID>356</GID>
<name>SEL_0</name></connection>
<intersection>-119.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211.5,-119.5,231.5,-119.5</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>231.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>226,-131.5,227.5,-131.5</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<connection>
<GID>359</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215,-129.5,227.5,-129.5</points>
<connection>
<GID>356</GID>
<name>IN_1</name></connection>
<connection>
<GID>360</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>206.5,-127.5,227.5,-127.5</points>
<connection>
<GID>356</GID>
<name>IN_2</name></connection>
<connection>
<GID>361</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>233.5,-128.5,252,-128.5</points>
<connection>
<GID>356</GID>
<name>OUT</name></connection>
<intersection>252 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>252,-128.5,252,-122.5</points>
<connection>
<GID>1050</GID>
<name>IN_0</name></connection>
<intersection>-128.5 1</intersection>
<intersection>-126 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>252,-126,294.5,-126</points>
<connection>
<GID>1200</GID>
<name>IN_0</name></connection>
<intersection>252 2</intersection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187,-136.5,187,-135.5</points>
<connection>
<GID>362</GID>
<name>SEL_1</name></connection>
<intersection>-135.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-135.5,187,-135.5</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188,-136.5,188,-132.5</points>
<connection>
<GID>362</GID>
<name>SEL_0</name></connection>
<intersection>-132.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-132.5,188,-132.5</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>188 0</intersection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>182.5,-144.5,184,-144.5</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<connection>
<GID>365</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>171.5,-142.5,184,-142.5</points>
<connection>
<GID>362</GID>
<name>IN_1</name></connection>
<connection>
<GID>366</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>163,-140.5,184,-140.5</points>
<connection>
<GID>362</GID>
<name>IN_2</name></connection>
<connection>
<GID>367</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-141.5,253.5,-141.5</points>
<connection>
<GID>362</GID>
<name>OUT</name></connection>
<intersection>253.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>253.5,-141.5,253.5,-135.5</points>
<connection>
<GID>1051</GID>
<name>IN_0</name></connection>
<intersection>-141.5 1</intersection>
<intersection>-140 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>253.5,-140,295,-140</points>
<connection>
<GID>1202</GID>
<name>IN_0</name></connection>
<intersection>253.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-149.5,231.5,-148.5</points>
<connection>
<GID>368</GID>
<name>SEL_1</name></connection>
<intersection>-148.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>212.5,-148.5,231.5,-148.5</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<intersection>231.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-149.5,232.5,-145.5</points>
<connection>
<GID>368</GID>
<name>SEL_0</name></connection>
<intersection>-145.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>212.5,-145.5,232.5,-145.5</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<intersection>232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-157.5,228.5,-157.5</points>
<connection>
<GID>368</GID>
<name>IN_0</name></connection>
<connection>
<GID>371</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216,-155.5,228.5,-155.5</points>
<connection>
<GID>368</GID>
<name>IN_1</name></connection>
<connection>
<GID>372</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>207.5,-153.5,228.5,-153.5</points>
<connection>
<GID>368</GID>
<name>IN_2</name></connection>
<connection>
<GID>373</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234.5,-154.5,252.5,-154.5</points>
<connection>
<GID>368</GID>
<name>OUT</name></connection>
<intersection>252.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>252.5,-154.5,252.5,-149</points>
<connection>
<GID>1052</GID>
<name>IN_0</name></connection>
<intersection>-154.5 1</intersection>
<intersection>-153 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>252.5,-153,295,-153</points>
<connection>
<GID>1204</GID>
<name>IN_0</name></connection>
<intersection>252.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-162.5,187.5,-161.5</points>
<connection>
<GID>374</GID>
<name>SEL_1</name></connection>
<intersection>-161.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,-161.5,187.5,-161.5</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-162.5,188.5,-158.5</points>
<connection>
<GID>374</GID>
<name>SEL_0</name></connection>
<intersection>-158.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,-158.5,188.5,-158.5</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>188.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>183,-170.5,184.5,-170.5</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<connection>
<GID>377</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-168.5,184.5,-168.5</points>
<connection>
<GID>374</GID>
<name>IN_1</name></connection>
<connection>
<GID>378</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>163.5,-166.5,184.5,-166.5</points>
<connection>
<GID>374</GID>
<name>IN_2</name></connection>
<connection>
<GID>379</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190.5,-167.5,252,-167.5</points>
<connection>
<GID>374</GID>
<name>OUT</name></connection>
<intersection>252 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>252,-167.5,252,-162</points>
<intersection>-167.5 1</intersection>
<intersection>-165.5 7</intersection>
<intersection>-162 10</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>252,-165.5,295,-165.5</points>
<connection>
<GID>1206</GID>
<name>IN_0</name></connection>
<intersection>252 2</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>252,-162,252.5,-162</points>
<connection>
<GID>1053</GID>
<name>IN_0</name></connection>
<intersection>252 2</intersection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233.5,-175.5,233.5,-174.5</points>
<connection>
<GID>380</GID>
<name>SEL_1</name></connection>
<intersection>-174.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>214,-174.5,233.5,-174.5</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>233.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234.5,-175.5,234.5,-171.5</points>
<connection>
<GID>380</GID>
<name>SEL_0</name></connection>
<intersection>-171.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>214,-171.5,234.5,-171.5</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>228.5,-183.5,230.5,-183.5</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<connection>
<GID>383</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217.5,-181.5,230.5,-181.5</points>
<connection>
<GID>380</GID>
<name>IN_1</name></connection>
<connection>
<GID>384</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>209,-179.5,230.5,-179.5</points>
<connection>
<GID>380</GID>
<name>IN_2</name></connection>
<connection>
<GID>385</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,-180.5,252,-180.5</points>
<connection>
<GID>380</GID>
<name>OUT</name></connection>
<intersection>252 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>252,-180.5,252,-175</points>
<connection>
<GID>1054</GID>
<name>IN_0</name></connection>
<intersection>-180.5 1</intersection>
<intersection>-179.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>252,-179.5,294.5,-179.5</points>
<connection>
<GID>1208</GID>
<name>IN_0</name></connection>
<intersection>252 2</intersection></hsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-189.5,188.5,-188.5</points>
<connection>
<GID>386</GID>
<name>SEL_1</name></connection>
<intersection>-188.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-188.5,188.5,-188.5</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>188.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,-189.5,189.5,-185.5</points>
<connection>
<GID>386</GID>
<name>SEL_0</name></connection>
<intersection>-185.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-185.5,189.5,-185.5</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>182.5,-197.5,185.5,-197.5</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<connection>
<GID>389</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>173,-195.5,185.5,-195.5</points>
<connection>
<GID>386</GID>
<name>IN_1</name></connection>
<connection>
<GID>390</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>164.5,-193.5,185.5,-193.5</points>
<connection>
<GID>386</GID>
<name>IN_2</name></connection>
<connection>
<GID>391</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>191.5,-194.5,252.5,-194.5</points>
<connection>
<GID>386</GID>
<name>OUT</name></connection>
<intersection>252.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>252.5,-194.5,252.5,-189</points>
<connection>
<GID>1055</GID>
<name>IN_0</name></connection>
<intersection>-194.5 1</intersection>
<intersection>-193.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>252.5,-193.5,294.5,-193.5</points>
<connection>
<GID>1210</GID>
<name>IN_0</name></connection>
<intersection>252.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233.5,-203.5,233.5,-202.5</points>
<connection>
<GID>392</GID>
<name>SEL_1</name></connection>
<intersection>-202.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>214.5,-202.5,233.5,-202.5</points>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<intersection>233.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234.5,-203.5,234.5,-199.5</points>
<connection>
<GID>392</GID>
<name>SEL_0</name></connection>
<intersection>-199.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>214.5,-199.5,234.5,-199.5</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>907</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>404,-63.5,404,-59</points>
<connection>
<GID>1133</GID>
<name>IN_0</name></connection>
<intersection>-63.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>404,-63.5,407.5,-63.5</points>
<connection>
<GID>1132</GID>
<name>IN_7</name></connection>
<intersection>404 0</intersection></hsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>229,-211.5,230.5,-211.5</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<connection>
<GID>395</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>908</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>403.5,-64.5,403.5,-56</points>
<intersection>-64.5 1</intersection>
<intersection>-56 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>403.5,-64.5,407.5,-64.5</points>
<connection>
<GID>1132</GID>
<name>IN_6</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>403.5,-56,405.5,-56</points>
<connection>
<GID>1134</GID>
<name>IN_0</name></connection>
<intersection>403.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-209.5,230.5,-209.5</points>
<connection>
<GID>392</GID>
<name>IN_1</name></connection>
<connection>
<GID>396</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>909</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>403,-65.5,403,-53</points>
<intersection>-65.5 1</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>403,-65.5,407.5,-65.5</points>
<connection>
<GID>1132</GID>
<name>IN_5</name></connection>
<intersection>403 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>403,-53,404,-53</points>
<connection>
<GID>1135</GID>
<name>IN_0</name></connection>
<intersection>403 0</intersection></hsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>209.5,-207.5,230.5,-207.5</points>
<connection>
<GID>392</GID>
<name>IN_2</name></connection>
<connection>
<GID>397</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>910</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>402.5,-66.5,402.5,-50</points>
<intersection>-66.5 1</intersection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>402.5,-66.5,407.5,-66.5</points>
<connection>
<GID>1132</GID>
<name>IN_4</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>402.5,-50,404,-50</points>
<connection>
<GID>1136</GID>
<name>IN_0</name></connection>
<intersection>402.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,-208.5,253,-208.5</points>
<connection>
<GID>392</GID>
<name>OUT</name></connection>
<intersection>253 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>253,-208.5,253,-203</points>
<connection>
<GID>1056</GID>
<name>IN_0</name></connection>
<intersection>-208.5 1</intersection>
<intersection>-206.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>253,-206.5,294,-206.5</points>
<connection>
<GID>1212</GID>
<name>IN_0</name></connection>
<intersection>253 2</intersection></hsegment></shape></wire>
<wire>
<ID>911</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>404,-75,404,-70.5</points>
<connection>
<GID>1140</GID>
<name>IN_0</name></connection>
<intersection>-70.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>404,-70.5,407.5,-70.5</points>
<connection>
<GID>1132</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-216.5,189,-215.5</points>
<connection>
<GID>398</GID>
<name>SEL_1</name></connection>
<intersection>-215.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170,-215.5,189,-215.5</points>
<connection>
<GID>399</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment></shape></wire>
<wire>
<ID>912</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>403.5,-78,403.5,-69.5</points>
<intersection>-78 2</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>403.5,-69.5,407.5,-69.5</points>
<connection>
<GID>1132</GID>
<name>IN_1</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>403.5,-78,404,-78</points>
<connection>
<GID>1139</GID>
<name>IN_0</name></connection>
<intersection>403.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,-216.5,190,-212.5</points>
<connection>
<GID>398</GID>
<name>SEL_0</name></connection>
<intersection>-212.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170,-212.5,190,-212.5</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<intersection>190 0</intersection></hsegment></shape></wire>
<wire>
<ID>913</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>403,-81,403,-68.5</points>
<intersection>-81 1</intersection>
<intersection>-68.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>403,-81,404,-81</points>
<connection>
<GID>1138</GID>
<name>IN_0</name></connection>
<intersection>403 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>403,-68.5,407.5,-68.5</points>
<connection>
<GID>1132</GID>
<name>IN_2</name></connection>
<intersection>403 0</intersection></hsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>184.5,-224.5,186,-224.5</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<connection>
<GID>401</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>914</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>402.5,-84,402.5,-67.5</points>
<intersection>-84 1</intersection>
<intersection>-67.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>402.5,-84,404,-84</points>
<connection>
<GID>1137</GID>
<name>IN_0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>402.5,-67.5,407.5,-67.5</points>
<connection>
<GID>1132</GID>
<name>IN_3</name></connection>
<intersection>402.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>173.5,-222.5,186,-222.5</points>
<connection>
<GID>398</GID>
<name>IN_1</name></connection>
<connection>
<GID>402</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>915</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380.5,-63,380.5,-58.5</points>
<connection>
<GID>1142</GID>
<name>IN_0</name></connection>
<intersection>-63 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>380.5,-63,384,-63</points>
<connection>
<GID>1141</GID>
<name>IN_7</name></connection>
<intersection>380.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-220.5,186,-220.5</points>
<connection>
<GID>398</GID>
<name>IN_2</name></connection>
<connection>
<GID>403</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>916</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380,-64,380,-55.5</points>
<intersection>-64 1</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380,-64,384,-64</points>
<connection>
<GID>1141</GID>
<name>IN_6</name></connection>
<intersection>380 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>380,-55.5,380.5,-55.5</points>
<connection>
<GID>1143</GID>
<name>IN_0</name></connection>
<intersection>380 0</intersection></hsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-221,252,-221</points>
<intersection>192 4</intersection>
<intersection>252 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>252,-221,252,-216</points>
<connection>
<GID>1057</GID>
<name>IN_0</name></connection>
<intersection>-221 1</intersection>
<intersection>-219 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>192,-221.5,192,-221</points>
<connection>
<GID>398</GID>
<name>OUT</name></connection>
<intersection>-221 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>252,-219,294,-219</points>
<connection>
<GID>1214</GID>
<name>IN_0</name></connection>
<intersection>252 2</intersection></hsegment></shape></wire>
<wire>
<ID>917</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379.5,-65,379.5,-52.5</points>
<intersection>-65 1</intersection>
<intersection>-52.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379.5,-65,384,-65</points>
<connection>
<GID>1141</GID>
<name>IN_5</name></connection>
<intersection>379.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>379.5,-52.5,380.5,-52.5</points>
<connection>
<GID>1144</GID>
<name>IN_0</name></connection>
<intersection>379.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237,-229.5,237,-228.5</points>
<connection>
<GID>404</GID>
<name>SEL_1</name></connection>
<intersection>-228.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>217,-228.5,237,-228.5</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>237 0</intersection></hsegment></shape></wire>
<wire>
<ID>918</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379,-66,379,-49.5</points>
<intersection>-66 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,-66,384,-66</points>
<connection>
<GID>1141</GID>
<name>IN_4</name></connection>
<intersection>379 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>379,-49.5,380.5,-49.5</points>
<connection>
<GID>1145</GID>
<name>IN_0</name></connection>
<intersection>379 0</intersection></hsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,-229.5,238,-225.5</points>
<connection>
<GID>404</GID>
<name>SEL_0</name></connection>
<intersection>-225.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>217,-225.5,238,-225.5</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment></shape></wire>
<wire>
<ID>919</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380.5,-74.5,380.5,-70</points>
<connection>
<GID>1149</GID>
<name>IN_0</name></connection>
<intersection>-70 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>380.5,-70,384,-70</points>
<connection>
<GID>1141</GID>
<name>IN_0</name></connection>
<intersection>380.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>231.5,-237.5,234,-237.5</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<connection>
<GID>407</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>920</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380,-77.5,380,-69</points>
<intersection>-77.5 2</intersection>
<intersection>-69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380,-69,384,-69</points>
<connection>
<GID>1141</GID>
<name>IN_1</name></connection>
<intersection>380 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>380,-77.5,380.5,-77.5</points>
<connection>
<GID>1148</GID>
<name>IN_0</name></connection>
<intersection>380 0</intersection></hsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220.5,-235.5,234,-235.5</points>
<connection>
<GID>404</GID>
<name>IN_1</name></connection>
<connection>
<GID>408</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>921</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379.5,-80.5,379.5,-68</points>
<intersection>-80.5 1</intersection>
<intersection>-68 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379.5,-80.5,380.5,-80.5</points>
<connection>
<GID>1147</GID>
<name>IN_0</name></connection>
<intersection>379.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>379.5,-68,384,-68</points>
<connection>
<GID>1141</GID>
<name>IN_2</name></connection>
<intersection>379.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212,-233.5,234,-233.5</points>
<connection>
<GID>404</GID>
<name>IN_2</name></connection>
<connection>
<GID>409</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>922</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379,-83.5,379,-67</points>
<intersection>-83.5 1</intersection>
<intersection>-67 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,-83.5,380.5,-83.5</points>
<connection>
<GID>1146</GID>
<name>IN_0</name></connection>
<intersection>379 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>379,-67,384,-67</points>
<connection>
<GID>1141</GID>
<name>IN_3</name></connection>
<intersection>379 0</intersection></hsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-234.5,252.5,-234.5</points>
<connection>
<GID>404</GID>
<name>OUT</name></connection>
<intersection>252.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>252.5,-234.5,252.5,-229</points>
<connection>
<GID>1058</GID>
<name>IN_0</name></connection>
<intersection>-234.5 1</intersection>
<intersection>-233 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>252.5,-233,294,-233</points>
<connection>
<GID>1216</GID>
<name>IN_0</name></connection>
<intersection>252.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,-243.5,189.5,-242.5</points>
<connection>
<GID>410</GID>
<name>SEL_1</name></connection>
<intersection>-242.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171,-242.5,189.5,-242.5</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,-243.5,190.5,-239.5</points>
<connection>
<GID>410</GID>
<name>SEL_0</name></connection>
<intersection>-239.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171,-239.5,190.5,-239.5</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>185.5,-251.5,186.5,-251.5</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<connection>
<GID>413</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174.5,-249.5,186.5,-249.5</points>
<connection>
<GID>410</GID>
<name>IN_1</name></connection>
<connection>
<GID>414</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166,-247.5,186.5,-247.5</points>
<connection>
<GID>410</GID>
<name>IN_2</name></connection>
<connection>
<GID>415</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192.5,-248.5,251.5,-248.5</points>
<connection>
<GID>410</GID>
<name>OUT</name></connection>
<intersection>251.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>251.5,-248.5,251.5,-242.5</points>
<connection>
<GID>1059</GID>
<name>IN_0</name></connection>
<intersection>-248.5 1</intersection>
<intersection>-247 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>251.5,-247,294.5,-247</points>
<connection>
<GID>1218</GID>
<name>IN_0</name></connection>
<intersection>251.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>232,-49.5,296,-49.5</points>
<intersection>232 6</intersection>
<intersection>248 2</intersection>
<intersection>296 5</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>248,-49.5,248,-46.5</points>
<connection>
<GID>1024</GID>
<name>IN_0</name></connection>
<intersection>-49.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>296,-51.5,296,-49.5</points>
<connection>
<GID>1186</GID>
<name>IN_0</name></connection>
<intersection>-49.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>232,-51.5,232,-49.5</points>
<connection>
<GID>246</GID>
<name>OUT</name></connection>
<intersection>-49.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-60,84.5,-55.5</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>-60 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>84.5,-60,88,-60</points>
<connection>
<GID>422</GID>
<name>IN_7</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-61,84,-52.5</points>
<intersection>-61 1</intersection>
<intersection>-52.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-61,88,-61</points>
<connection>
<GID>422</GID>
<name>IN_6</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84,-52.5,84.5,-52.5</points>
<connection>
<GID>426</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-62,83.5,-49.5</points>
<intersection>-62 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-62,88,-62</points>
<connection>
<GID>422</GID>
<name>IN_5</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,-49.5,84.5,-49.5</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-63,83,-46.5</points>
<intersection>-63 1</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-63,88,-63</points>
<connection>
<GID>422</GID>
<name>IN_4</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83,-46.5,84.5,-46.5</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-71.5,84.5,-67</points>
<connection>
<GID>434</GID>
<name>IN_0</name></connection>
<intersection>-67 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>84.5,-67,88,-67</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-74.5,84,-66</points>
<intersection>-74.5 2</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-66,88,-66</points>
<connection>
<GID>422</GID>
<name>IN_1</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84,-74.5,84.5,-74.5</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-77.5,83.5,-65</points>
<intersection>-77.5 1</intersection>
<intersection>-65 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-77.5,84.5,-77.5</points>
<connection>
<GID>432</GID>
<name>IN_0</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,-65,88,-65</points>
<connection>
<GID>422</GID>
<name>IN_2</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-80.5,83,-64</points>
<intersection>-80.5 1</intersection>
<intersection>-64 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-80.5,84.5,-80.5</points>
<connection>
<GID>431</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83,-64,88,-64</points>
<connection>
<GID>422</GID>
<name>IN_3</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-60,63.5,-55.5</points>
<connection>
<GID>445</GID>
<name>IN_0</name></connection>
<intersection>-60 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>63.5,-60,67,-60</points>
<connection>
<GID>444</GID>
<name>IN_7</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-61,63,-52.5</points>
<intersection>-61 1</intersection>
<intersection>-52.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-61,67,-61</points>
<connection>
<GID>444</GID>
<name>IN_6</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-52.5,63.5,-52.5</points>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-62,62.5,-49.5</points>
<intersection>-62 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-62,67,-62</points>
<connection>
<GID>444</GID>
<name>IN_5</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-49.5,63.5,-49.5</points>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>953</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>302,-51.5,306,-51.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<connection>
<GID>1186</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-63,62,-46.5</points>
<intersection>-63 1</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-63,67,-63</points>
<connection>
<GID>444</GID>
<name>IN_4</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62,-46.5,63.5,-46.5</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>954</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>291.5,-53.5,296,-53.5</points>
<connection>
<GID>1186</GID>
<name>clock</name></connection>
<connection>
<GID>1187</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-71.5,63.5,-67</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<intersection>-67 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>63.5,-67,67,-67</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>955</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292,-65.5,296.5,-65.5</points>
<connection>
<GID>1190</GID>
<name>clock</name></connection>
<connection>
<GID>1189</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-74.5,63,-66</points>
<intersection>-74.5 2</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-66,67,-66</points>
<connection>
<GID>444</GID>
<name>IN_1</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-74.5,63.5,-74.5</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>956</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,-64.5,304,-63.5</points>
<intersection>-64.5 1</intersection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-64.5,306,-64.5</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>304 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>302.5,-63.5,304,-63.5</points>
<connection>
<GID>1190</GID>
<name>OUT_0</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-77.5,62.5,-65</points>
<intersection>-77.5 1</intersection>
<intersection>-65 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-77.5,63.5,-77.5</points>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-65,67,-65</points>
<connection>
<GID>444</GID>
<name>IN_2</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>957</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-78,294.5,-78</points>
<connection>
<GID>1192</GID>
<name>clock</name></connection>
<connection>
<GID>1191</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-80.5,62,-64</points>
<intersection>-80.5 1</intersection>
<intersection>-64 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-80.5,63.5,-80.5</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62,-64,67,-64</points>
<connection>
<GID>444</GID>
<name>IN_3</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>958</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,-77.5,303.5,-76</points>
<intersection>-77.5 2</intersection>
<intersection>-76 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>300.5,-76,303.5,-76</points>
<connection>
<GID>1192</GID>
<name>OUT_0</name></connection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-77.5,307,-77.5</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>959</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290.5,-91,294.5,-91</points>
<connection>
<GID>1193</GID>
<name>IN_0</name></connection>
<intersection>294.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>294.5,-91.5,294.5,-91</points>
<connection>
<GID>1194</GID>
<name>clock</name></connection>
<intersection>-91 1</intersection></vsegment></shape></wire>
<wire>
<ID>960</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,-90.5,303.5,-89.5</points>
<intersection>-90.5 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-90.5,307,-90.5</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300.5,-89.5,303.5,-89.5</points>
<connection>
<GID>1194</GID>
<name>OUT_0</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>961</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290.5,-103.5,295,-103.5</points>
<connection>
<GID>1196</GID>
<name>clock</name></connection>
<connection>
<GID>1195</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>962</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,-103.5,304,-101.5</points>
<intersection>-103.5 1</intersection>
<intersection>-101.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-103.5,307,-103.5</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>304 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,-101.5,304,-101.5</points>
<connection>
<GID>1196</GID>
<name>OUT_0</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>963</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-115.5,294.5,-115.5</points>
<connection>
<GID>1198</GID>
<name>clock</name></connection>
<connection>
<GID>1197</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>964</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,-115.5,303.5,-113.5</points>
<intersection>-115.5 1</intersection>
<intersection>-113.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-115.5,307,-115.5</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300.5,-113.5,303.5,-113.5</points>
<connection>
<GID>1198</GID>
<name>OUT_0</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>186.527,63.765,1964.53,-853.235</PageViewport>
<gate>
<ID>416</ID>
<type>DA_FROM</type>
<position>357,-140</position>
<input>
<ID>IN_0</ID>213 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_MUX_OUT</lparam></gate>
<gate>
<ID>417</ID>
<type>DA_FROM</type>
<position>357,-143</position>
<input>
<ID>IN_0</ID>214 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B2_IN</lparam></gate>
<gate>
<ID>418</ID>
<type>DE_TO</type>
<position>390,-139</position>
<input>
<ID>IN_0</ID>241 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_ULA</lparam></gate>
<gate>
<ID>419</ID>
<type>DE_TO</type>
<position>385,-148</position>
<input>
<ID>IN_0</ID>242 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B3_IN</lparam></gate>
<gate>
<ID>421</ID>
<type>AI_XOR2</type>
<position>379.5,-169.5</position>
<input>
<ID>IN_0</ID>352 </input>
<input>
<ID>IN_1</ID>243 </input>
<output>
<ID>OUT</ID>249 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>423</ID>
<type>AI_XOR2</type>
<position>371.5,-170.5</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>252 </input>
<output>
<ID>OUT</ID>243 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>425</ID>
<type>AE_OR3</type>
<position>379.5,-177.5</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>247 </input>
<input>
<ID>IN_2</ID>244 </input>
<output>
<ID>OUT</ID>364 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>427</ID>
<type>AA_AND2</type>
<position>371,-175.5</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>252 </input>
<output>
<ID>OUT</ID>248 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>429</ID>
<type>AA_AND2</type>
<position>371.5,-181</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>253 </input>
<output>
<ID>OUT</ID>247 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>435</ID>
<type>AA_AND2</type>
<position>371.5,-186</position>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>351 </input>
<output>
<ID>OUT</ID>244 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>436</ID>
<type>AA_MUX_2x1</type>
<position>385.5,-168.5</position>
<input>
<ID>IN_0</ID>249 </input>
<input>
<ID>IN_1</ID>354 </input>
<output>
<ID>OUT</ID>355 </output>
<input>
<ID>SEL_0</ID>353 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>437</ID>
<type>AE_SMALL_INVERTER</type>
<position>366,-182</position>
<input>
<ID>IN_0</ID>352 </input>
<output>
<ID>OUT_0</ID>253 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>438</ID>
<type>AE_SMALL_INVERTER</type>
<position>366,-187</position>
<input>
<ID>IN_0</ID>352 </input>
<output>
<ID>OUT_0</ID>351 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>439</ID>
<type>DA_FROM</type>
<position>357,-160.5</position>
<input>
<ID>IN_0</ID>353 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>440</ID>
<type>DA_FROM</type>
<position>357,-163.5</position>
<input>
<ID>IN_0</ID>354 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_SOMA</lparam></gate>
<gate>
<ID>441</ID>
<type>DA_FROM</type>
<position>357,-166.5</position>
<input>
<ID>IN_0</ID>352 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_ACC_OUT</lparam></gate>
<gate>
<ID>442</ID>
<type>DA_FROM</type>
<position>357.5,-169.5</position>
<input>
<ID>IN_0</ID>251 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_MUX_OUT</lparam></gate>
<gate>
<ID>443</ID>
<type>DA_FROM</type>
<position>357.5,-172.5</position>
<input>
<ID>IN_0</ID>252 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B3_IN</lparam></gate>
<gate>
<ID>453</ID>
<type>DE_TO</type>
<position>391.5,-168.5</position>
<input>
<ID>IN_0</ID>355 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_ULA</lparam></gate>
<gate>
<ID>455</ID>
<type>DE_TO</type>
<position>385.5,-177.5</position>
<input>
<ID>IN_0</ID>364 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B4_IN</lparam></gate>
<gate>
<ID>456</ID>
<type>DE_TO</type>
<position>292,-132.5</position>
<input>
<ID>IN_0</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_SOMA</lparam></gate>
<gate>
<ID>458</ID>
<type>DE_TO</type>
<position>292,-135.5</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_SOMA</lparam></gate>
<gate>
<ID>459</ID>
<type>DA_FROM</type>
<position>430,-140</position>
<input>
<ID>IN_0</ID>371 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_MUX_OUT</lparam></gate>
<gate>
<ID>461</ID>
<type>DA_FROM</type>
<position>430,-143</position>
<input>
<ID>IN_0</ID>384 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B10_IN</lparam></gate>
<gate>
<ID>462</ID>
<type>DE_TO</type>
<position>463,-139</position>
<input>
<ID>IN_0</ID>390 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_ULA</lparam></gate>
<gate>
<ID>463</ID>
<type>DE_TO</type>
<position>458,-148</position>
<input>
<ID>IN_0</ID>391 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B11_IN</lparam></gate>
<gate>
<ID>464</ID>
<type>AI_XOR2</type>
<position>452.5,-169.5</position>
<input>
<ID>IN_0</ID>402 </input>
<input>
<ID>IN_1</ID>392 </input>
<output>
<ID>OUT</ID>397 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>465</ID>
<type>AI_XOR2</type>
<position>444.5,-170.5</position>
<input>
<ID>IN_0</ID>398 </input>
<input>
<ID>IN_1</ID>399 </input>
<output>
<ID>OUT</ID>392 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>466</ID>
<type>AE_OR3</type>
<position>452.5,-177.5</position>
<input>
<ID>IN_0</ID>395 </input>
<input>
<ID>IN_1</ID>394 </input>
<input>
<ID>IN_2</ID>393 </input>
<output>
<ID>OUT</ID>406 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>467</ID>
<type>AA_AND2</type>
<position>444.5,-175.5</position>
<input>
<ID>IN_0</ID>398 </input>
<input>
<ID>IN_1</ID>399 </input>
<output>
<ID>OUT</ID>395 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>468</ID>
<type>AA_AND2</type>
<position>444.5,-181</position>
<input>
<ID>IN_0</ID>398 </input>
<input>
<ID>IN_1</ID>400 </input>
<output>
<ID>OUT</ID>394 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>469</ID>
<type>AA_AND2</type>
<position>444.5,-186</position>
<input>
<ID>IN_0</ID>399 </input>
<input>
<ID>IN_1</ID>401 </input>
<output>
<ID>OUT</ID>393 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>470</ID>
<type>AA_MUX_2x1</type>
<position>458.5,-168.5</position>
<input>
<ID>IN_0</ID>397 </input>
<input>
<ID>IN_1</ID>404 </input>
<output>
<ID>OUT</ID>405 </output>
<input>
<ID>SEL_0</ID>403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>471</ID>
<type>AE_SMALL_INVERTER</type>
<position>439,-182</position>
<input>
<ID>IN_0</ID>402 </input>
<output>
<ID>OUT_0</ID>400 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>472</ID>
<type>AE_SMALL_INVERTER</type>
<position>439,-187</position>
<input>
<ID>IN_0</ID>402 </input>
<output>
<ID>OUT_0</ID>401 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>473</ID>
<type>DA_FROM</type>
<position>430,-160.5</position>
<input>
<ID>IN_0</ID>403 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>474</ID>
<type>DA_FROM</type>
<position>430,-163.5</position>
<input>
<ID>IN_0</ID>404 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_SOMA</lparam></gate>
<gate>
<ID>475</ID>
<type>DA_FROM</type>
<position>430,-166.5</position>
<input>
<ID>IN_0</ID>402 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_ACC_OUT</lparam></gate>
<gate>
<ID>476</ID>
<type>DA_FROM</type>
<position>430.5,-169.5</position>
<input>
<ID>IN_0</ID>398 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_MUX_OUT</lparam></gate>
<gate>
<ID>477</ID>
<type>DA_FROM</type>
<position>430.5,-172.5</position>
<input>
<ID>IN_0</ID>399 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B11_IN</lparam></gate>
<gate>
<ID>478</ID>
<type>DE_TO</type>
<position>464,-168.5</position>
<input>
<ID>IN_0</ID>405 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_ULA</lparam></gate>
<gate>
<ID>868</ID>
<type>AA_LABEL</type>
<position>289.5,-96.5</position>
<gparam>LABEL_TEXT Sinais de Controle</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>479</ID>
<type>DE_TO</type>
<position>458.5,-177.5</position>
<input>
<ID>IN_0</ID>406 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B12_IN</lparam></gate>
<gate>
<ID>869</ID>
<type>AA_LABEL</type>
<position>270.5,-106</position>
<gparam>LABEL_TEXT OP_ULA</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>480</ID>
<type>DE_TO</type>
<position>292,-138.5</position>
<input>
<ID>IN_0</ID>154 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_SOMA</lparam></gate>
<gate>
<ID>482</ID>
<type>AI_XOR2</type>
<position>452,-140</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>370 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>483</ID>
<type>DE_TO</type>
<position>292,-141.5</position>
<input>
<ID>IN_0</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_SOMA</lparam></gate>
<gate>
<ID>484</ID>
<type>AI_XOR2</type>
<position>444,-141</position>
<input>
<ID>IN_0</ID>371 </input>
<input>
<ID>IN_1</ID>384 </input>
<output>
<ID>OUT</ID>366 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>485</ID>
<type>AE_OR3</type>
<position>452,-148</position>
<input>
<ID>IN_0</ID>369 </input>
<input>
<ID>IN_1</ID>368 </input>
<input>
<ID>IN_2</ID>367 </input>
<output>
<ID>OUT</ID>391 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>486</ID>
<type>DE_TO</type>
<position>292,-159.5</position>
<input>
<ID>IN_0</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_SOMA</lparam></gate>
<gate>
<ID>487</ID>
<type>AA_AND2</type>
<position>444,-146</position>
<input>
<ID>IN_0</ID>371 </input>
<input>
<ID>IN_1</ID>384 </input>
<output>
<ID>OUT</ID>369 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>488</ID>
<type>AA_AND2</type>
<position>444,-151.5</position>
<input>
<ID>IN_0</ID>371 </input>
<input>
<ID>IN_1</ID>385 </input>
<output>
<ID>OUT</ID>368 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>489</ID>
<type>AA_AND2</type>
<position>444,-156.5</position>
<input>
<ID>IN_0</ID>384 </input>
<input>
<ID>IN_1</ID>386 </input>
<output>
<ID>OUT</ID>367 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>490</ID>
<type>AA_MUX_2x1</type>
<position>458,-139</position>
<input>
<ID>IN_0</ID>370 </input>
<input>
<ID>IN_1</ID>389 </input>
<output>
<ID>OUT</ID>390 </output>
<input>
<ID>SEL_0</ID>388 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>491</ID>
<type>AE_SMALL_INVERTER</type>
<position>438.5,-152.5</position>
<input>
<ID>IN_0</ID>387 </input>
<output>
<ID>OUT_0</ID>385 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>492</ID>
<type>AE_SMALL_INVERTER</type>
<position>438.5,-157.5</position>
<input>
<ID>IN_0</ID>387 </input>
<output>
<ID>OUT_0</ID>386 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>493</ID>
<type>DA_FROM</type>
<position>429.5,-131</position>
<input>
<ID>IN_0</ID>388 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>494</ID>
<type>DE_TO</type>
<position>384,-90.5</position>
<input>
<ID>IN_0</ID>396 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BO_IN</lparam></gate>
<gate>
<ID>495</ID>
<type>DA_FROM</type>
<position>429.5,-134</position>
<input>
<ID>IN_0</ID>389 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_SOMA</lparam></gate>
<gate>
<ID>496</ID>
<type>FF_GND</type>
<position>381,-92.5</position>
<output>
<ID>OUT_0</ID>396 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>497</ID>
<type>DA_FROM</type>
<position>429.5,-137</position>
<input>
<ID>IN_0</ID>387 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_ACC_OUT</lparam></gate>
<gate>
<ID>498</ID>
<type>AI_XOR2</type>
<position>451,-78.5</position>
<input>
<ID>IN_0</ID>426 </input>
<input>
<ID>IN_1</ID>408 </input>
<output>
<ID>OUT</ID>417 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>499</ID>
<type>AI_XOR2</type>
<position>443,-79.5</position>
<input>
<ID>IN_0</ID>418 </input>
<input>
<ID>IN_1</ID>420 </input>
<output>
<ID>OUT</ID>408 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>500</ID>
<type>AE_OR3</type>
<position>451,-86.5</position>
<input>
<ID>IN_0</ID>411 </input>
<input>
<ID>IN_1</ID>410 </input>
<input>
<ID>IN_2</ID>409 </input>
<output>
<ID>OUT</ID>435 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>501</ID>
<type>AA_AND2</type>
<position>443,-84.5</position>
<input>
<ID>IN_0</ID>418 </input>
<input>
<ID>IN_1</ID>420 </input>
<output>
<ID>OUT</ID>411 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>502</ID>
<type>AA_AND2</type>
<position>443,-90</position>
<input>
<ID>IN_0</ID>418 </input>
<input>
<ID>IN_1</ID>424 </input>
<output>
<ID>OUT</ID>410 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>503</ID>
<type>AA_AND2</type>
<position>443,-95</position>
<input>
<ID>IN_0</ID>420 </input>
<input>
<ID>IN_1</ID>425 </input>
<output>
<ID>OUT</ID>409 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>504</ID>
<type>AA_MUX_2x1</type>
<position>457,-77.5</position>
<input>
<ID>IN_0</ID>417 </input>
<input>
<ID>IN_1</ID>428 </input>
<output>
<ID>OUT</ID>430 </output>
<input>
<ID>SEL_0</ID>427 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>505</ID>
<type>AE_SMALL_INVERTER</type>
<position>437.5,-91</position>
<input>
<ID>IN_0</ID>426 </input>
<output>
<ID>OUT_0</ID>424 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>506</ID>
<type>AE_SMALL_INVERTER</type>
<position>437.5,-96</position>
<input>
<ID>IN_0</ID>426 </input>
<output>
<ID>OUT_0</ID>425 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>507</ID>
<type>DA_FROM</type>
<position>428.5,-69.5</position>
<input>
<ID>IN_0</ID>427 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>508</ID>
<type>DA_FROM</type>
<position>428.5,-72.5</position>
<input>
<ID>IN_0</ID>428 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_SOMA</lparam></gate>
<gate>
<ID>509</ID>
<type>DA_FROM</type>
<position>428.5,-75.5</position>
<input>
<ID>IN_0</ID>426 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_ACC_OUT</lparam></gate>
<gate>
<ID>510</ID>
<type>DA_FROM</type>
<position>429,-78.5</position>
<input>
<ID>IN_0</ID>418 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_MUX_OUT</lparam></gate>
<gate>
<ID>511</ID>
<type>DA_FROM</type>
<position>429,-81.5</position>
<input>
<ID>IN_0</ID>420 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B8_IN</lparam></gate>
<gate>
<ID>512</ID>
<type>DE_TO</type>
<position>462,-77.5</position>
<input>
<ID>IN_0</ID>430 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_ULA</lparam></gate>
<gate>
<ID>513</ID>
<type>DE_TO</type>
<position>457,-86.5</position>
<input>
<ID>IN_0</ID>435 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B9_IN</lparam></gate>
<gate>
<ID>514</ID>
<type>AI_XOR2</type>
<position>451.5,-108</position>
<input>
<ID>IN_0</ID>459 </input>
<input>
<ID>IN_1</ID>450 </input>
<output>
<ID>OUT</ID>454 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>515</ID>
<type>AI_XOR2</type>
<position>443.5,-109</position>
<input>
<ID>IN_0</ID>455 </input>
<input>
<ID>IN_1</ID>456 </input>
<output>
<ID>OUT</ID>450 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>516</ID>
<type>AA_LABEL</type>
<position>377.5,-44.5</position>
<gparam>LABEL_TEXT Unidade Logica e Aritmetica - ULA</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>517</ID>
<type>AE_OR3</type>
<position>451.5,-116</position>
<input>
<ID>IN_0</ID>453 </input>
<input>
<ID>IN_1</ID>452 </input>
<input>
<ID>IN_2</ID>451 </input>
<output>
<ID>OUT</ID>463 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>518</ID>
<type>AI_XOR2</type>
<position>378,-78.5</position>
<input>
<ID>IN_0</ID>429 </input>
<input>
<ID>IN_1</ID>412 </input>
<output>
<ID>OUT</ID>416 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>519</ID>
<type>AI_XOR2</type>
<position>370,-79.5</position>
<input>
<ID>IN_0</ID>419 </input>
<input>
<ID>IN_1</ID>421 </input>
<output>
<ID>OUT</ID>412 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>520</ID>
<type>AE_OR3</type>
<position>378,-86.5</position>
<input>
<ID>IN_0</ID>415 </input>
<input>
<ID>IN_1</ID>414 </input>
<input>
<ID>IN_2</ID>413 </input>
<output>
<ID>OUT</ID>434 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>521</ID>
<type>AA_AND2</type>
<position>370,-84.5</position>
<input>
<ID>IN_0</ID>419 </input>
<input>
<ID>IN_1</ID>421 </input>
<output>
<ID>OUT</ID>415 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>522</ID>
<type>AA_AND2</type>
<position>370,-90</position>
<input>
<ID>IN_0</ID>419 </input>
<input>
<ID>IN_1</ID>422 </input>
<output>
<ID>OUT</ID>414 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>523</ID>
<type>AA_AND2</type>
<position>370,-95</position>
<input>
<ID>IN_0</ID>421 </input>
<input>
<ID>IN_1</ID>423 </input>
<output>
<ID>OUT</ID>413 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>524</ID>
<type>AA_MUX_2x1</type>
<position>384,-77.5</position>
<input>
<ID>IN_0</ID>416 </input>
<input>
<ID>IN_1</ID>432 </input>
<output>
<ID>OUT</ID>433 </output>
<input>
<ID>SEL_0</ID>431 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>525</ID>
<type>AA_AND2</type>
<position>443.5,-114</position>
<input>
<ID>IN_0</ID>455 </input>
<input>
<ID>IN_1</ID>456 </input>
<output>
<ID>OUT</ID>453 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>526</ID>
<type>AA_AND2</type>
<position>443.5,-119.5</position>
<input>
<ID>IN_0</ID>455 </input>
<input>
<ID>IN_1</ID>457 </input>
<output>
<ID>OUT</ID>452 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>527</ID>
<type>AA_AND2</type>
<position>443.5,-124.5</position>
<input>
<ID>IN_0</ID>456 </input>
<input>
<ID>IN_1</ID>458 </input>
<output>
<ID>OUT</ID>451 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>528</ID>
<type>AA_MUX_2x1</type>
<position>457.5,-107</position>
<input>
<ID>IN_0</ID>454 </input>
<input>
<ID>IN_1</ID>461 </input>
<output>
<ID>OUT</ID>462 </output>
<input>
<ID>SEL_0</ID>460 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>529</ID>
<type>AE_SMALL_INVERTER</type>
<position>438,-120.5</position>
<input>
<ID>IN_0</ID>459 </input>
<output>
<ID>OUT_0</ID>457 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>530</ID>
<type>AE_SMALL_INVERTER</type>
<position>364.5,-91</position>
<input>
<ID>IN_0</ID>429 </input>
<output>
<ID>OUT_0</ID>422 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>531</ID>
<type>AE_SMALL_INVERTER</type>
<position>364.5,-96</position>
<input>
<ID>IN_0</ID>429 </input>
<output>
<ID>OUT_0</ID>423 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>532</ID>
<type>AE_SMALL_INVERTER</type>
<position>438,-125.5</position>
<input>
<ID>IN_0</ID>459 </input>
<output>
<ID>OUT_0</ID>458 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>533</ID>
<type>DA_FROM</type>
<position>429,-99</position>
<input>
<ID>IN_0</ID>460 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>534</ID>
<type>DA_FROM</type>
<position>429,-102</position>
<input>
<ID>IN_0</ID>461 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_SOMA</lparam></gate>
<gate>
<ID>535</ID>
<type>DA_FROM</type>
<position>429,-105</position>
<input>
<ID>IN_0</ID>459 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_ACC_OUT</lparam></gate>
<gate>
<ID>536</ID>
<type>DA_FROM</type>
<position>429.5,-108</position>
<input>
<ID>IN_0</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_MUX_OUT</lparam></gate>
<gate>
<ID>537</ID>
<type>DA_FROM</type>
<position>429.5,-111</position>
<input>
<ID>IN_0</ID>456 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B9_IN</lparam></gate>
<gate>
<ID>538</ID>
<type>DE_TO</type>
<position>463,-107</position>
<input>
<ID>IN_0</ID>462 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_ULA</lparam></gate>
<gate>
<ID>149</ID>
<type>AE_FULLADDER_4BIT</type>
<position>283,-136</position>
<input>
<ID>IN_0</ID>365 </input>
<input>
<ID>IN_1</ID>380 </input>
<input>
<ID>IN_2</ID>381 </input>
<input>
<ID>IN_3</ID>382 </input>
<input>
<ID>IN_B_0</ID>203 </input>
<input>
<ID>IN_B_1</ID>202 </input>
<input>
<ID>IN_B_2</ID>201 </input>
<input>
<ID>IN_B_3</ID>157 </input>
<output>
<ID>OUT_0</ID>156 </output>
<output>
<ID>OUT_1</ID>153 </output>
<output>
<ID>OUT_2</ID>154 </output>
<output>
<ID>OUT_3</ID>155 </output>
<input>
<ID>carry_in</ID>613 </input>
<output>
<ID>carry_out</ID>610 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>539</ID>
<type>DE_TO</type>
<position>457.5,-116</position>
<input>
<ID>IN_0</ID>463 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B10_IN</lparam></gate>
<gate>
<ID>540</ID>
<type>DA_FROM</type>
<position>358.5,-266.5</position>
<input>
<ID>IN_0</ID>470 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_MUX_OUT</lparam></gate>
<gate>
<ID>541</ID>
<type>DA_FROM</type>
<position>358.5,-269.5</position>
<input>
<ID>IN_0</ID>471 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B6_IN</lparam></gate>
<gate>
<ID>152</ID>
<type>DA_FROM</type>
<position>272,-134</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_ACC_OUT</lparam></gate>
<gate>
<ID>542</ID>
<type>DE_TO</type>
<position>391.5,-265.5</position>
<input>
<ID>IN_0</ID>477 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_ULA</lparam></gate>
<gate>
<ID>543</ID>
<type>DE_TO</type>
<position>386.5,-274.5</position>
<input>
<ID>IN_0</ID>478 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B7_IN</lparam></gate>
<gate>
<ID>544</ID>
<type>AI_XOR2</type>
<position>381,-296</position>
<input>
<ID>IN_0</ID>488 </input>
<input>
<ID>IN_1</ID>479 </input>
<output>
<ID>OUT</ID>483 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>545</ID>
<type>AI_XOR2</type>
<position>373,-297</position>
<input>
<ID>IN_0</ID>484 </input>
<input>
<ID>IN_1</ID>485 </input>
<output>
<ID>OUT</ID>479 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>546</ID>
<type>AE_OR3</type>
<position>381,-304</position>
<input>
<ID>IN_0</ID>482 </input>
<input>
<ID>IN_1</ID>481 </input>
<input>
<ID>IN_2</ID>480 </input>
<output>
<ID>OUT</ID>492 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>547</ID>
<type>AA_AND2</type>
<position>373,-302.5</position>
<input>
<ID>IN_0</ID>484 </input>
<input>
<ID>IN_1</ID>485 </input>
<output>
<ID>OUT</ID>482 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>158</ID>
<type>DA_FROM</type>
<position>272,-138</position>
<input>
<ID>IN_0</ID>365 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_MUX_OUT</lparam></gate>
<gate>
<ID>548</ID>
<type>AA_AND2</type>
<position>373,-307.5</position>
<input>
<ID>IN_0</ID>484 </input>
<input>
<ID>IN_1</ID>486 </input>
<output>
<ID>OUT</ID>481 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>549</ID>
<type>AA_AND2</type>
<position>373,-312.5</position>
<input>
<ID>IN_0</ID>485 </input>
<input>
<ID>IN_1</ID>487 </input>
<output>
<ID>OUT</ID>480 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>550</ID>
<type>AA_MUX_2x1</type>
<position>387,-295</position>
<input>
<ID>IN_0</ID>483 </input>
<input>
<ID>IN_1</ID>490 </input>
<output>
<ID>OUT</ID>491 </output>
<input>
<ID>SEL_0</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>551</ID>
<type>AE_SMALL_INVERTER</type>
<position>367.5,-308.5</position>
<input>
<ID>IN_0</ID>488 </input>
<output>
<ID>OUT_0</ID>486 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>552</ID>
<type>AE_SMALL_INVERTER</type>
<position>367.5,-313.5</position>
<input>
<ID>IN_0</ID>488 </input>
<output>
<ID>OUT_0</ID>487 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>553</ID>
<type>DA_FROM</type>
<position>355.5,-69.5</position>
<input>
<ID>IN_0</ID>431 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>554</ID>
<type>DA_FROM</type>
<position>358.5,-287</position>
<input>
<ID>IN_0</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>555</ID>
<type>DA_FROM</type>
<position>355.5,-72.5</position>
<input>
<ID>IN_0</ID>432 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_SOMA</lparam></gate>
<gate>
<ID>556</ID>
<type>DA_FROM</type>
<position>355.5,-75.5</position>
<input>
<ID>IN_0</ID>429 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_ACC_OUT</lparam></gate>
<gate>
<ID>557</ID>
<type>DA_FROM</type>
<position>356,-78.5</position>
<input>
<ID>IN_0</ID>419 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_MUX_OUT</lparam></gate>
<gate>
<ID>558</ID>
<type>DA_FROM</type>
<position>356,-81.5</position>
<input>
<ID>IN_0</ID>421 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BO_IN</lparam></gate>
<gate>
<ID>559</ID>
<type>DE_TO</type>
<position>389,-77.5</position>
<input>
<ID>IN_0</ID>433 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_ULA</lparam></gate>
<gate>
<ID>560</ID>
<type>DE_TO</type>
<position>384,-86.5</position>
<input>
<ID>IN_0</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B1_IN</lparam></gate>
<gate>
<ID>561</ID>
<type>DA_FROM</type>
<position>358.5,-290</position>
<input>
<ID>IN_0</ID>490 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_SOMA</lparam></gate>
<gate>
<ID>562</ID>
<type>DA_FROM</type>
<position>358.5,-293</position>
<input>
<ID>IN_0</ID>488 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_ACC_OUT</lparam></gate>
<gate>
<ID>563</ID>
<type>AI_XOR2</type>
<position>378.5,-108</position>
<input>
<ID>IN_0</ID>445 </input>
<input>
<ID>IN_1</ID>436 </input>
<output>
<ID>OUT</ID>440 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>564</ID>
<type>AI_XOR2</type>
<position>370.5,-109</position>
<input>
<ID>IN_0</ID>441 </input>
<input>
<ID>IN_1</ID>442 </input>
<output>
<ID>OUT</ID>436 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>565</ID>
<type>AE_OR3</type>
<position>378.5,-116</position>
<input>
<ID>IN_0</ID>439 </input>
<input>
<ID>IN_1</ID>438 </input>
<input>
<ID>IN_2</ID>437 </input>
<output>
<ID>OUT</ID>449 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>566</ID>
<type>AA_AND2</type>
<position>370.5,-114</position>
<input>
<ID>IN_0</ID>441 </input>
<input>
<ID>IN_1</ID>442 </input>
<output>
<ID>OUT</ID>439 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>567</ID>
<type>AA_AND2</type>
<position>370.5,-119.5</position>
<input>
<ID>IN_0</ID>441 </input>
<input>
<ID>IN_1</ID>443 </input>
<output>
<ID>OUT</ID>438 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>568</ID>
<type>AA_AND2</type>
<position>370.5,-124.5</position>
<input>
<ID>IN_0</ID>442 </input>
<input>
<ID>IN_1</ID>444 </input>
<output>
<ID>OUT</ID>437 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>569</ID>
<type>AA_MUX_2x1</type>
<position>384.5,-107</position>
<input>
<ID>IN_0</ID>440 </input>
<input>
<ID>IN_1</ID>447 </input>
<output>
<ID>OUT</ID>448 </output>
<input>
<ID>SEL_0</ID>446 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>570</ID>
<type>AE_SMALL_INVERTER</type>
<position>365,-120.5</position>
<input>
<ID>IN_0</ID>445 </input>
<output>
<ID>OUT_0</ID>443 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>571</ID>
<type>AE_SMALL_INVERTER</type>
<position>365,-125.5</position>
<input>
<ID>IN_0</ID>445 </input>
<output>
<ID>OUT_0</ID>444 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>572</ID>
<type>DA_FROM</type>
<position>356,-99</position>
<input>
<ID>IN_0</ID>446 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>573</ID>
<type>DA_FROM</type>
<position>356,-102</position>
<input>
<ID>IN_0</ID>447 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_SOMA</lparam></gate>
<gate>
<ID>574</ID>
<type>DA_FROM</type>
<position>356,-105</position>
<input>
<ID>IN_0</ID>445 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_ACC_OUT</lparam></gate>
<gate>
<ID>575</ID>
<type>DA_FROM</type>
<position>356.5,-108</position>
<input>
<ID>IN_0</ID>441 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_MUX_OUT</lparam></gate>
<gate>
<ID>576</ID>
<type>DA_FROM</type>
<position>356.5,-111</position>
<input>
<ID>IN_0</ID>442 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B1_IN</lparam></gate>
<gate>
<ID>187</ID>
<type>DA_FROM</type>
<position>272,-141.5</position>
<input>
<ID>IN_0</ID>380 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_MUX_OUT</lparam></gate>
<gate>
<ID>577</ID>
<type>DE_TO</type>
<position>390,-107</position>
<input>
<ID>IN_0</ID>448 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_ULA</lparam></gate>
<gate>
<ID>578</ID>
<type>DE_TO</type>
<position>384.5,-116</position>
<input>
<ID>IN_0</ID>449 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B2_IN</lparam></gate>
<gate>
<ID>579</ID>
<type>DA_FROM</type>
<position>359,-296</position>
<input>
<ID>IN_0</ID>484 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_MUX_OUT</lparam></gate>
<gate>
<ID>581</ID>
<type>DA_FROM</type>
<position>359,-299</position>
<input>
<ID>IN_0</ID>485 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B7_IN</lparam></gate>
<gate>
<ID>583</ID>
<type>DE_TO</type>
<position>392.5,-295</position>
<input>
<ID>IN_0</ID>491 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_ULA</lparam></gate>
<gate>
<ID>585</ID>
<type>DE_TO</type>
<position>387,-304</position>
<input>
<ID>IN_0</ID>492 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B8_IN</lparam></gate>
<gate>
<ID>587</ID>
<type>DA_FROM</type>
<position>431.5,-266.5</position>
<input>
<ID>IN_0</ID>499 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_MUX_OUT</lparam></gate>
<gate>
<ID>589</ID>
<type>DA_FROM</type>
<position>431.5,-269.5</position>
<input>
<ID>IN_0</ID>500 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B14_IN</lparam></gate>
<gate>
<ID>591</ID>
<type>DE_TO</type>
<position>464.5,-265.5</position>
<input>
<ID>IN_0</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_ULA</lparam></gate>
<gate>
<ID>593</ID>
<type>DE_TO</type>
<position>459.5,-274.5</position>
<input>
<ID>IN_0</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B15_IN</lparam></gate>
<gate>
<ID>594</ID>
<type>AI_XOR2</type>
<position>454,-296</position>
<input>
<ID>IN_0</ID>518 </input>
<input>
<ID>IN_1</ID>508 </input>
<output>
<ID>OUT</ID>513 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>DA_FROM</type>
<position>272,-144.5</position>
<input>
<ID>IN_0</ID>381 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_MUX_OUT</lparam></gate>
<gate>
<ID>595</ID>
<type>AI_XOR2</type>
<position>446,-297</position>
<input>
<ID>IN_0</ID>514 </input>
<input>
<ID>IN_1</ID>515 </input>
<output>
<ID>OUT</ID>508 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>596</ID>
<type>AE_OR3</type>
<position>454,-304</position>
<input>
<ID>IN_0</ID>511 </input>
<input>
<ID>IN_1</ID>510 </input>
<input>
<ID>IN_2</ID>509 </input>
<output>
<ID>OUT</ID>580 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>597</ID>
<type>AA_AND2</type>
<position>446,-302.5</position>
<input>
<ID>IN_0</ID>514 </input>
<input>
<ID>IN_1</ID>515 </input>
<output>
<ID>OUT</ID>511 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>598</ID>
<type>AA_AND2</type>
<position>446,-307.5</position>
<input>
<ID>IN_0</ID>514 </input>
<input>
<ID>IN_1</ID>516 </input>
<output>
<ID>OUT</ID>510 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>599</ID>
<type>AA_AND2</type>
<position>446,-312.5</position>
<input>
<ID>IN_0</ID>515 </input>
<input>
<ID>IN_1</ID>517 </input>
<output>
<ID>OUT</ID>509 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>600</ID>
<type>AA_MUX_2x1</type>
<position>460,-295</position>
<input>
<ID>IN_0</ID>513 </input>
<input>
<ID>IN_1</ID>520 </input>
<output>
<ID>OUT</ID>521 </output>
<input>
<ID>SEL_0</ID>519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>601</ID>
<type>AE_SMALL_INVERTER</type>
<position>440.5,-308.5</position>
<input>
<ID>IN_0</ID>518 </input>
<output>
<ID>OUT_0</ID>516 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>602</ID>
<type>AE_SMALL_INVERTER</type>
<position>440.5,-313.5</position>
<input>
<ID>IN_0</ID>518 </input>
<output>
<ID>OUT_0</ID>517 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>603</ID>
<type>DA_FROM</type>
<position>431.5,-287</position>
<input>
<ID>IN_0</ID>519 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>604</ID>
<type>DA_FROM</type>
<position>431.5,-290</position>
<input>
<ID>IN_0</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_SOMA</lparam></gate>
<gate>
<ID>605</ID>
<type>DA_FROM</type>
<position>431.5,-293</position>
<input>
<ID>IN_0</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_ACC_OUT</lparam></gate>
<gate>
<ID>606</ID>
<type>DA_FROM</type>
<position>432,-296</position>
<input>
<ID>IN_0</ID>514 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_MUX_OUT</lparam></gate>
<gate>
<ID>607</ID>
<type>DA_FROM</type>
<position>432,-299</position>
<input>
<ID>IN_0</ID>515 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B15_IN</lparam></gate>
<gate>
<ID>608</ID>
<type>DE_TO</type>
<position>465.5,-295</position>
<input>
<ID>IN_0</ID>521 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_ULA</lparam></gate>
<gate>
<ID>609</ID>
<type>DE_TO</type>
<position>292,-162.5</position>
<input>
<ID>IN_0</ID>383 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_SOMA</lparam></gate>
<gate>
<ID>610</ID>
<type>DE_TO</type>
<position>292,-165.5</position>
<input>
<ID>IN_0</ID>407 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_SOMA</lparam></gate>
<gate>
<ID>611</ID>
<type>DE_TO</type>
<position>292,-168.5</position>
<input>
<ID>IN_0</ID>464 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_SOMA</lparam></gate>
<gate>
<ID>612</ID>
<type>AI_XOR2</type>
<position>453.5,-266.5</position>
<input>
<ID>IN_0</ID>503 </input>
<input>
<ID>IN_1</ID>494 </input>
<output>
<ID>OUT</ID>498 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>613</ID>
<type>AE_FULLADDER_4BIT</type>
<position>283,-163</position>
<input>
<ID>IN_0</ID>582 </input>
<input>
<ID>IN_1</ID>583 </input>
<input>
<ID>IN_2</ID>584 </input>
<input>
<ID>IN_3</ID>585 </input>
<input>
<ID>IN_B_0</ID>581 </input>
<input>
<ID>IN_B_1</ID>523 </input>
<input>
<ID>IN_B_2</ID>522 </input>
<input>
<ID>IN_B_3</ID>512 </input>
<output>
<ID>OUT_0</ID>493 </output>
<output>
<ID>OUT_1</ID>383 </output>
<output>
<ID>OUT_2</ID>407 </output>
<output>
<ID>OUT_3</ID>464 </output>
<input>
<ID>carry_in</ID>610 </input>
<output>
<ID>carry_out</ID>611 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>614</ID>
<type>AI_XOR2</type>
<position>445.5,-267.5</position>
<input>
<ID>IN_0</ID>499 </input>
<input>
<ID>IN_1</ID>500 </input>
<output>
<ID>OUT</ID>494 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>615</ID>
<type>AE_OR3</type>
<position>453.5,-274.5</position>
<input>
<ID>IN_0</ID>497 </input>
<input>
<ID>IN_1</ID>496 </input>
<input>
<ID>IN_2</ID>495 </input>
<output>
<ID>OUT</ID>507 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>616</ID>
<type>DA_FROM</type>
<position>272,-161</position>
<input>
<ID>IN_0</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_ACC_OUT</lparam></gate>
<gate>
<ID>617</ID>
<type>AA_AND2</type>
<position>445.5,-272.5</position>
<input>
<ID>IN_0</ID>499 </input>
<input>
<ID>IN_1</ID>500 </input>
<output>
<ID>OUT</ID>497 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>618</ID>
<type>AA_AND2</type>
<position>445.5,-278</position>
<input>
<ID>IN_0</ID>499 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>496 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>619</ID>
<type>AA_AND2</type>
<position>445.5,-283</position>
<input>
<ID>IN_0</ID>500 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>495 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>620</ID>
<type>AA_MUX_2x1</type>
<position>459.5,-265.5</position>
<input>
<ID>IN_0</ID>498 </input>
<input>
<ID>IN_1</ID>505 </input>
<output>
<ID>OUT</ID>506 </output>
<input>
<ID>SEL_0</ID>504 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>621</ID>
<type>AE_SMALL_INVERTER</type>
<position>440,-279</position>
<input>
<ID>IN_0</ID>503 </input>
<output>
<ID>OUT_0</ID>501 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>622</ID>
<type>AE_SMALL_INVERTER</type>
<position>440,-284</position>
<input>
<ID>IN_0</ID>503 </input>
<output>
<ID>OUT_0</ID>502 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>623</ID>
<type>DA_FROM</type>
<position>272,-165</position>
<input>
<ID>IN_0</ID>582 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_MUX_OUT</lparam></gate>
<gate>
<ID>624</ID>
<type>DA_FROM</type>
<position>431,-257.5</position>
<input>
<ID>IN_0</ID>504 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>625</ID>
<type>DA_FROM</type>
<position>272,-168.5</position>
<input>
<ID>IN_0</ID>583 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_MUX_OUT</lparam></gate>
<gate>
<ID>626</ID>
<type>AI_XOR2</type>
<position>380.5,-266.5</position>
<input>
<ID>IN_0</ID>474 </input>
<input>
<ID>IN_1</ID>465 </input>
<output>
<ID>OUT</ID>469 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>627</ID>
<type>DA_FROM</type>
<position>272,-171.5</position>
<input>
<ID>IN_0</ID>584 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_MUX_OUT</lparam></gate>
<gate>
<ID>628</ID>
<type>DA_FROM</type>
<position>431,-260.5</position>
<input>
<ID>IN_0</ID>505 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_SOMA</lparam></gate>
<gate>
<ID>629</ID>
<type>AI_XOR2</type>
<position>372.5,-267.5</position>
<input>
<ID>IN_0</ID>470 </input>
<input>
<ID>IN_1</ID>471 </input>
<output>
<ID>OUT</ID>465 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>630</ID>
<type>AE_OR3</type>
<position>380.5,-274.5</position>
<input>
<ID>IN_0</ID>468 </input>
<input>
<ID>IN_1</ID>467 </input>
<input>
<ID>IN_2</ID>466 </input>
<output>
<ID>OUT</ID>478 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>631</ID>
<type>DA_FROM</type>
<position>272,-174.5</position>
<input>
<ID>IN_0</ID>585 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_MUX_OUT</lparam></gate>
<gate>
<ID>632</ID>
<type>DA_FROM</type>
<position>431,-263.5</position>
<input>
<ID>IN_0</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_ACC_OUT</lparam></gate>
<gate>
<ID>633</ID>
<type>AI_XOR2</type>
<position>452.5,-205</position>
<input>
<ID>IN_0</ID>542 </input>
<input>
<ID>IN_1</ID>524 </input>
<output>
<ID>OUT</ID>533 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>634</ID>
<type>AI_XOR2</type>
<position>444.5,-206</position>
<input>
<ID>IN_0</ID>534 </input>
<input>
<ID>IN_1</ID>536 </input>
<output>
<ID>OUT</ID>524 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>635</ID>
<type>AE_OR3</type>
<position>452.5,-213</position>
<input>
<ID>IN_0</ID>527 </input>
<input>
<ID>IN_1</ID>526 </input>
<input>
<ID>IN_2</ID>525 </input>
<output>
<ID>OUT</ID>551 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>636</ID>
<type>AA_AND2</type>
<position>444.5,-211</position>
<input>
<ID>IN_0</ID>534 </input>
<input>
<ID>IN_1</ID>536 </input>
<output>
<ID>OUT</ID>527 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>637</ID>
<type>AA_AND2</type>
<position>444.5,-216.5</position>
<input>
<ID>IN_0</ID>534 </input>
<input>
<ID>IN_1</ID>540 </input>
<output>
<ID>OUT</ID>526 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>638</ID>
<type>AA_AND2</type>
<position>372,-272.5</position>
<input>
<ID>IN_0</ID>470 </input>
<input>
<ID>IN_1</ID>471 </input>
<output>
<ID>OUT</ID>468 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>639</ID>
<type>AA_AND2</type>
<position>444.5,-221.5</position>
<input>
<ID>IN_0</ID>536 </input>
<input>
<ID>IN_1</ID>541 </input>
<output>
<ID>OUT</ID>525 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>640</ID>
<type>AA_MUX_2x1</type>
<position>458.5,-204</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>544 </input>
<output>
<ID>OUT</ID>546 </output>
<input>
<ID>SEL_0</ID>543 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>641</ID>
<type>AE_SMALL_INVERTER</type>
<position>439,-217.5</position>
<input>
<ID>IN_0</ID>542 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>642</ID>
<type>AE_SMALL_INVERTER</type>
<position>439,-222.5</position>
<input>
<ID>IN_0</ID>542 </input>
<output>
<ID>OUT_0</ID>541 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>643</ID>
<type>AA_AND2</type>
<position>372.5,-278</position>
<input>
<ID>IN_0</ID>470 </input>
<input>
<ID>IN_1</ID>472 </input>
<output>
<ID>OUT</ID>467 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>644</ID>
<type>DA_FROM</type>
<position>430,-196</position>
<input>
<ID>IN_0</ID>543 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>645</ID>
<type>AA_AND2</type>
<position>372.5,-283</position>
<input>
<ID>IN_0</ID>471 </input>
<input>
<ID>IN_1</ID>473 </input>
<output>
<ID>OUT</ID>466 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>646</ID>
<type>DA_FROM</type>
<position>430,-199</position>
<input>
<ID>IN_0</ID>544 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_SOMA</lparam></gate>
<gate>
<ID>647</ID>
<type>AA_MUX_2x1</type>
<position>386.5,-265.5</position>
<input>
<ID>IN_0</ID>469 </input>
<input>
<ID>IN_1</ID>476 </input>
<output>
<ID>OUT</ID>477 </output>
<input>
<ID>SEL_0</ID>475 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>648</ID>
<type>DA_FROM</type>
<position>430,-202</position>
<input>
<ID>IN_0</ID>542 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_ACC_OUT</lparam></gate>
<gate>
<ID>649</ID>
<type>AE_SMALL_INVERTER</type>
<position>367,-279</position>
<input>
<ID>IN_0</ID>474 </input>
<output>
<ID>OUT_0</ID>472 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>650</ID>
<type>DA_FROM</type>
<position>430.5,-205</position>
<input>
<ID>IN_0</ID>534 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_MUX_OUT</lparam></gate>
<gate>
<ID>261</ID>
<type>AA_LABEL</type>
<position>356,-26</position>
<gparam>LABEL_TEXT Prof.  Angelo Zanini / Nuncio Perrella</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>651</ID>
<type>DA_FROM</type>
<position>430.5,-208</position>
<input>
<ID>IN_0</ID>536 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B12_IN</lparam></gate>
<gate>
<ID>652</ID>
<type>AE_SMALL_INVERTER</type>
<position>367,-284</position>
<input>
<ID>IN_0</ID>474 </input>
<output>
<ID>OUT_0</ID>473 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>653</ID>
<type>DE_TO</type>
<position>463.5,-204</position>
<input>
<ID>IN_0</ID>546 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_ULA</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_LABEL</type>
<position>364.5,-15</position>
<gparam>LABEL_TEXT PROCESSADOR BIP IMT - MAUA 2022</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>654</ID>
<type>DE_TO</type>
<position>458.5,-213</position>
<input>
<ID>IN_0</ID>551 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B13_IN</lparam></gate>
<gate>
<ID>655</ID>
<type>DA_FROM</type>
<position>358,-257.5</position>
<input>
<ID>IN_0</ID>475 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>656</ID>
<type>AI_XOR2</type>
<position>453,-234.5</position>
<input>
<ID>IN_0</ID>575 </input>
<input>
<ID>IN_1</ID>566 </input>
<output>
<ID>OUT</ID>570 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>657</ID>
<type>AI_XOR2</type>
<position>445,-235.5</position>
<input>
<ID>IN_0</ID>571 </input>
<input>
<ID>IN_1</ID>572 </input>
<output>
<ID>OUT</ID>566 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>658</ID>
<type>DA_FROM</type>
<position>358,-260.5</position>
<input>
<ID>IN_0</ID>476 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_SOMA</lparam></gate>
<gate>
<ID>659</ID>
<type>AE_OR3</type>
<position>453,-242.5</position>
<input>
<ID>IN_0</ID>569 </input>
<input>
<ID>IN_1</ID>568 </input>
<input>
<ID>IN_2</ID>567 </input>
<output>
<ID>OUT</ID>579 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>660</ID>
<type>DA_FROM</type>
<position>358,-263.5</position>
<input>
<ID>IN_0</ID>474 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_ACC_OUT</lparam></gate>
<gate>
<ID>661</ID>
<type>AI_XOR2</type>
<position>379.5,-205</position>
<input>
<ID>IN_0</ID>545 </input>
<input>
<ID>IN_1</ID>528 </input>
<output>
<ID>OUT</ID>532 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>662</ID>
<type>AI_XOR2</type>
<position>371.5,-206</position>
<input>
<ID>IN_0</ID>535 </input>
<input>
<ID>IN_1</ID>537 </input>
<output>
<ID>OUT</ID>528 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>663</ID>
<type>AE_OR3</type>
<position>379.5,-213</position>
<input>
<ID>IN_0</ID>531 </input>
<input>
<ID>IN_1</ID>530 </input>
<input>
<ID>IN_2</ID>529 </input>
<output>
<ID>OUT</ID>550 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>664</ID>
<type>AA_AND2</type>
<position>371.5,-211</position>
<input>
<ID>IN_0</ID>535 </input>
<input>
<ID>IN_1</ID>537 </input>
<output>
<ID>OUT</ID>531 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>665</ID>
<type>AA_AND2</type>
<position>371.5,-216.5</position>
<input>
<ID>IN_0</ID>535 </input>
<input>
<ID>IN_1</ID>538 </input>
<output>
<ID>OUT</ID>530 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>666</ID>
<type>AA_AND2</type>
<position>371.5,-221.5</position>
<input>
<ID>IN_0</ID>537 </input>
<input>
<ID>IN_1</ID>539 </input>
<output>
<ID>OUT</ID>529 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>667</ID>
<type>AA_MUX_2x1</type>
<position>385.5,-204</position>
<input>
<ID>IN_0</ID>532 </input>
<input>
<ID>IN_1</ID>548 </input>
<output>
<ID>OUT</ID>549 </output>
<input>
<ID>SEL_0</ID>547 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>668</ID>
<type>AA_AND2</type>
<position>445,-240.5</position>
<input>
<ID>IN_0</ID>571 </input>
<input>
<ID>IN_1</ID>572 </input>
<output>
<ID>OUT</ID>569 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>DA_FROM</type>
<position>272,-147</position>
<input>
<ID>IN_0</ID>382 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_MUX_OUT</lparam></gate>
<gate>
<ID>669</ID>
<type>AA_AND2</type>
<position>445,-246</position>
<input>
<ID>IN_0</ID>571 </input>
<input>
<ID>IN_1</ID>573 </input>
<output>
<ID>OUT</ID>568 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>670</ID>
<type>AA_AND2</type>
<position>445,-251</position>
<input>
<ID>IN_0</ID>572 </input>
<input>
<ID>IN_1</ID>574 </input>
<output>
<ID>OUT</ID>567 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>671</ID>
<type>AA_MUX_2x1</type>
<position>459,-233.5</position>
<input>
<ID>IN_0</ID>570 </input>
<input>
<ID>IN_1</ID>577 </input>
<output>
<ID>OUT</ID>578 </output>
<input>
<ID>SEL_0</ID>576 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>672</ID>
<type>AE_SMALL_INVERTER</type>
<position>439.5,-247</position>
<input>
<ID>IN_0</ID>575 </input>
<output>
<ID>OUT_0</ID>573 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>673</ID>
<type>AE_SMALL_INVERTER</type>
<position>366,-217.5</position>
<input>
<ID>IN_0</ID>545 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>674</ID>
<type>AE_SMALL_INVERTER</type>
<position>366,-222.5</position>
<input>
<ID>IN_0</ID>545 </input>
<output>
<ID>OUT_0</ID>539 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>675</ID>
<type>AE_SMALL_INVERTER</type>
<position>439.5,-252</position>
<input>
<ID>IN_0</ID>575 </input>
<output>
<ID>OUT_0</ID>574 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>676</ID>
<type>DA_FROM</type>
<position>430.5,-225.5</position>
<input>
<ID>IN_0</ID>576 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>677</ID>
<type>DA_FROM</type>
<position>430.5,-228.5</position>
<input>
<ID>IN_0</ID>577 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_SOMA</lparam></gate>
<gate>
<ID>678</ID>
<type>DA_FROM</type>
<position>430.5,-231.5</position>
<input>
<ID>IN_0</ID>575 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_ACC_OUT</lparam></gate>
<gate>
<ID>679</ID>
<type>DA_FROM</type>
<position>431,-234.5</position>
<input>
<ID>IN_0</ID>571 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_MUX_OUT</lparam></gate>
<gate>
<ID>680</ID>
<type>DA_FROM</type>
<position>431,-237.5</position>
<input>
<ID>IN_0</ID>572 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B13_IN</lparam></gate>
<gate>
<ID>681</ID>
<type>DE_TO</type>
<position>464.5,-233.5</position>
<input>
<ID>IN_0</ID>578 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_ULA</lparam></gate>
<gate>
<ID>682</ID>
<type>DE_TO</type>
<position>459,-242.5</position>
<input>
<ID>IN_0</ID>579 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B14_IN</lparam></gate>
<gate>
<ID>683</ID>
<type>DA_FROM</type>
<position>357,-196</position>
<input>
<ID>IN_0</ID>547 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>684</ID>
<type>DA_FROM</type>
<position>357,-199</position>
<input>
<ID>IN_0</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_SOMA</lparam></gate>
<gate>
<ID>685</ID>
<type>DA_FROM</type>
<position>357,-202</position>
<input>
<ID>IN_0</ID>545 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_ACC_OUT</lparam></gate>
<gate>
<ID>296</ID>
<type>DA_FROM</type>
<position>272,-130.5</position>
<input>
<ID>IN_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_ACC_OUT</lparam></gate>
<gate>
<ID>686</ID>
<type>DA_FROM</type>
<position>357.5,-205</position>
<input>
<ID>IN_0</ID>535 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_MUX_OUT</lparam></gate>
<gate>
<ID>687</ID>
<type>DA_FROM</type>
<position>357.5,-208</position>
<input>
<ID>IN_0</ID>537 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B4_IN</lparam></gate>
<gate>
<ID>298</ID>
<type>DA_FROM</type>
<position>272,-127.5</position>
<input>
<ID>IN_0</ID>202 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_ACC_OUT</lparam></gate>
<gate>
<ID>688</ID>
<type>DE_TO</type>
<position>390.5,-204</position>
<input>
<ID>IN_0</ID>549 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_ULA</lparam></gate>
<gate>
<ID>689</ID>
<type>DE_TO</type>
<position>385.5,-213</position>
<input>
<ID>IN_0</ID>550 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B5_IN</lparam></gate>
<gate>
<ID>300</ID>
<type>DA_FROM</type>
<position>272,-124.5</position>
<input>
<ID>IN_0</ID>203 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_ACC_OUT</lparam></gate>
<gate>
<ID>690</ID>
<type>AI_XOR2</type>
<position>380,-234.5</position>
<input>
<ID>IN_0</ID>561 </input>
<input>
<ID>IN_1</ID>552 </input>
<output>
<ID>OUT</ID>556 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>301</ID>
<type>AI_XOR2</type>
<position>379,-140</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>204 </input>
<output>
<ID>OUT</ID>211 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>691</ID>
<type>AI_XOR2</type>
<position>372,-235.5</position>
<input>
<ID>IN_0</ID>557 </input>
<input>
<ID>IN_1</ID>558 </input>
<output>
<ID>OUT</ID>552 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>302</ID>
<type>AI_XOR2</type>
<position>371,-141</position>
<input>
<ID>IN_0</ID>213 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>692</ID>
<type>AE_OR3</type>
<position>380,-242.5</position>
<input>
<ID>IN_0</ID>555 </input>
<input>
<ID>IN_1</ID>554 </input>
<input>
<ID>IN_2</ID>553 </input>
<output>
<ID>OUT</ID>565 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>303</ID>
<type>AE_OR3</type>
<position>379,-148</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>206 </input>
<input>
<ID>IN_2</ID>205 </input>
<output>
<ID>OUT</ID>242 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>693</ID>
<type>AA_AND2</type>
<position>372,-240.5</position>
<input>
<ID>IN_0</ID>557 </input>
<input>
<ID>IN_1</ID>558 </input>
<output>
<ID>OUT</ID>555 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>694</ID>
<type>AA_AND2</type>
<position>372,-246</position>
<input>
<ID>IN_0</ID>557 </input>
<input>
<ID>IN_1</ID>559 </input>
<output>
<ID>OUT</ID>554 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>695</ID>
<type>AA_AND2</type>
<position>372,-251</position>
<input>
<ID>IN_0</ID>558 </input>
<input>
<ID>IN_1</ID>560 </input>
<output>
<ID>OUT</ID>553 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>696</ID>
<type>AA_MUX_2x1</type>
<position>386,-233.5</position>
<input>
<ID>IN_0</ID>556 </input>
<input>
<ID>IN_1</ID>563 </input>
<output>
<ID>OUT</ID>564 </output>
<input>
<ID>SEL_0</ID>562 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>697</ID>
<type>AE_SMALL_INVERTER</type>
<position>366.5,-247</position>
<input>
<ID>IN_0</ID>561 </input>
<output>
<ID>OUT_0</ID>559 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>698</ID>
<type>AE_SMALL_INVERTER</type>
<position>366.5,-252</position>
<input>
<ID>IN_0</ID>561 </input>
<output>
<ID>OUT_0</ID>560 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>309</ID>
<type>AA_AND2</type>
<position>371,-146</position>
<input>
<ID>IN_0</ID>213 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>699</ID>
<type>DA_FROM</type>
<position>357.5,-225.5</position>
<input>
<ID>IN_0</ID>562 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>700</ID>
<type>DA_FROM</type>
<position>357.5,-228.5</position>
<input>
<ID>IN_0</ID>563 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_SOMA</lparam></gate>
<gate>
<ID>701</ID>
<type>DA_FROM</type>
<position>357.5,-231.5</position>
<input>
<ID>IN_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_ACC_OUT</lparam></gate>
<gate>
<ID>702</ID>
<type>DA_FROM</type>
<position>358,-234.5</position>
<input>
<ID>IN_0</ID>557 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_MUX_OUT</lparam></gate>
<gate>
<ID>313</ID>
<type>AA_AND2</type>
<position>371,-151.5</position>
<input>
<ID>IN_0</ID>213 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>703</ID>
<type>DA_FROM</type>
<position>358,-237.5</position>
<input>
<ID>IN_0</ID>558 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B5_IN</lparam></gate>
<gate>
<ID>314</ID>
<type>AA_AND2</type>
<position>371,-156.5</position>
<input>
<ID>IN_0</ID>214 </input>
<input>
<ID>IN_1</ID>216 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>704</ID>
<type>DE_TO</type>
<position>391.5,-233.5</position>
<input>
<ID>IN_0</ID>564 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_ULA</lparam></gate>
<gate>
<ID>315</ID>
<type>AA_MUX_2x1</type>
<position>385,-139</position>
<input>
<ID>IN_0</ID>211 </input>
<input>
<ID>IN_1</ID>238 </input>
<output>
<ID>OUT</ID>241 </output>
<input>
<ID>SEL_0</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>705</ID>
<type>DE_TO</type>
<position>386,-242.5</position>
<input>
<ID>IN_0</ID>565 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B6_IN</lparam></gate>
<gate>
<ID>316</ID>
<type>AE_SMALL_INVERTER</type>
<position>365.5,-152.5</position>
<input>
<ID>IN_0</ID>218 </input>
<output>
<ID>OUT_0</ID>215 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>706</ID>
<type>DA_FROM</type>
<position>272,-157.5</position>
<input>
<ID>IN_0</ID>522 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_ACC_OUT</lparam></gate>
<gate>
<ID>707</ID>
<type>GA_LED</type>
<position>468,-304</position>
<input>
<ID>N_in0</ID>580 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>318</ID>
<type>AE_SMALL_INVERTER</type>
<position>365.5,-157.5</position>
<input>
<ID>IN_0</ID>218 </input>
<output>
<ID>OUT_0</ID>216 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>708</ID>
<type>DA_FROM</type>
<position>272,-154.5</position>
<input>
<ID>IN_0</ID>523 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_ACC_OUT</lparam></gate>
<gate>
<ID>320</ID>
<type>DA_FROM</type>
<position>356.5,-131</position>
<input>
<ID>IN_0</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>709</ID>
<type>DA_FROM</type>
<position>272,-151.5</position>
<input>
<ID>IN_0</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_ACC_OUT</lparam></gate>
<gate>
<ID>710</ID>
<type>DE_TO</type>
<position>292,-186.5</position>
<input>
<ID>IN_0</ID>589 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_SOMA</lparam></gate>
<gate>
<ID>322</ID>
<type>DA_FROM</type>
<position>356.5,-134</position>
<input>
<ID>IN_0</ID>238 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_SOMA</lparam></gate>
<gate>
<ID>711</ID>
<type>DE_TO</type>
<position>292,-189.5</position>
<input>
<ID>IN_0</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_SOMA</lparam></gate>
<gate>
<ID>712</ID>
<type>DE_TO</type>
<position>292,-192.5</position>
<input>
<ID>IN_0</ID>587 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_SOMA</lparam></gate>
<gate>
<ID>324</ID>
<type>DA_FROM</type>
<position>356.5,-137</position>
<input>
<ID>IN_0</ID>218 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_ACC_OUT</lparam></gate>
<gate>
<ID>713</ID>
<type>DE_TO</type>
<position>292,-195.5</position>
<input>
<ID>IN_0</ID>588 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_SOMA</lparam></gate>
<gate>
<ID>714</ID>
<type>AE_FULLADDER_4BIT</type>
<position>283,-190</position>
<input>
<ID>IN_0</ID>594 </input>
<input>
<ID>IN_1</ID>595 </input>
<input>
<ID>IN_2</ID>596 </input>
<input>
<ID>IN_3</ID>597 </input>
<input>
<ID>IN_B_0</ID>593 </input>
<input>
<ID>IN_B_1</ID>592 </input>
<input>
<ID>IN_B_2</ID>591 </input>
<input>
<ID>IN_B_3</ID>590 </input>
<output>
<ID>OUT_0</ID>589 </output>
<output>
<ID>OUT_1</ID>586 </output>
<output>
<ID>OUT_2</ID>587 </output>
<output>
<ID>OUT_3</ID>588 </output>
<input>
<ID>carry_in</ID>611 </input>
<output>
<ID>carry_out</ID>612 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>715</ID>
<type>DA_FROM</type>
<position>272,-188</position>
<input>
<ID>IN_0</ID>590 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_ACC_OUT</lparam></gate>
<gate>
<ID>716</ID>
<type>DA_FROM</type>
<position>272,-192</position>
<input>
<ID>IN_0</ID>594 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_MUX_OUT</lparam></gate>
<gate>
<ID>717</ID>
<type>DA_FROM</type>
<position>272,-195.5</position>
<input>
<ID>IN_0</ID>595 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_MUX_OUT</lparam></gate>
<gate>
<ID>718</ID>
<type>DA_FROM</type>
<position>272,-198.5</position>
<input>
<ID>IN_0</ID>596 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_MUX_OUT</lparam></gate>
<gate>
<ID>719</ID>
<type>DA_FROM</type>
<position>272,-201.5</position>
<input>
<ID>IN_0</ID>597 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_MUX_OUT</lparam></gate>
<gate>
<ID>720</ID>
<type>DA_FROM</type>
<position>272,-184.5</position>
<input>
<ID>IN_0</ID>591 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_ACC_OUT</lparam></gate>
<gate>
<ID>721</ID>
<type>DA_FROM</type>
<position>272.5,-181.5</position>
<input>
<ID>IN_0</ID>592 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_ACC_OUT</lparam></gate>
<gate>
<ID>722</ID>
<type>DA_FROM</type>
<position>272,-178.5</position>
<input>
<ID>IN_0</ID>593 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_ACC_OUT</lparam></gate>
<gate>
<ID>723</ID>
<type>DE_TO</type>
<position>292,-213.5</position>
<input>
<ID>IN_0</ID>601 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_SOMA</lparam></gate>
<gate>
<ID>724</ID>
<type>DE_TO</type>
<position>292,-216.5</position>
<input>
<ID>IN_0</ID>598 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_SOMA</lparam></gate>
<gate>
<ID>725</ID>
<type>DE_TO</type>
<position>292,-219.5</position>
<input>
<ID>IN_0</ID>599 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_SOMA</lparam></gate>
<gate>
<ID>726</ID>
<type>DE_TO</type>
<position>292,-222.5</position>
<input>
<ID>IN_0</ID>600 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_SOMA</lparam></gate>
<gate>
<ID>727</ID>
<type>AE_FULLADDER_4BIT</type>
<position>283,-217</position>
<input>
<ID>IN_0</ID>606 </input>
<input>
<ID>IN_1</ID>607 </input>
<input>
<ID>IN_2</ID>608 </input>
<input>
<ID>IN_3</ID>609 </input>
<input>
<ID>IN_B_0</ID>605 </input>
<input>
<ID>IN_B_1</ID>604 </input>
<input>
<ID>IN_B_2</ID>603 </input>
<input>
<ID>IN_B_3</ID>602 </input>
<output>
<ID>OUT_0</ID>601 </output>
<output>
<ID>OUT_1</ID>598 </output>
<output>
<ID>OUT_2</ID>599 </output>
<output>
<ID>OUT_3</ID>600 </output>
<input>
<ID>carry_in</ID>612 </input>
<output>
<ID>carry_out</ID>614 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>728</ID>
<type>DA_FROM</type>
<position>272,-215</position>
<input>
<ID>IN_0</ID>602 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_ACC_OUT</lparam></gate>
<gate>
<ID>729</ID>
<type>DA_FROM</type>
<position>272,-219</position>
<input>
<ID>IN_0</ID>606 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_MUX_OUT</lparam></gate>
<gate>
<ID>730</ID>
<type>DA_FROM</type>
<position>272,-222.5</position>
<input>
<ID>IN_0</ID>607 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_MUX_OUT</lparam></gate>
<gate>
<ID>731</ID>
<type>DA_FROM</type>
<position>272,-225.5</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_MUX_OUT</lparam></gate>
<gate>
<ID>732</ID>
<type>DA_FROM</type>
<position>272,-228.5</position>
<input>
<ID>IN_0</ID>609 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_MUX_OUT</lparam></gate>
<gate>
<ID>733</ID>
<type>DA_FROM</type>
<position>272,-211.5</position>
<input>
<ID>IN_0</ID>603 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_ACC_OUT</lparam></gate>
<gate>
<ID>734</ID>
<type>DA_FROM</type>
<position>272,-208.5</position>
<input>
<ID>IN_0</ID>604 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_ACC_OUT</lparam></gate>
<gate>
<ID>735</ID>
<type>DA_FROM</type>
<position>272,-205.5</position>
<input>
<ID>IN_0</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_ACC_OUT</lparam></gate>
<gate>
<ID>737</ID>
<type>FF_GND</type>
<position>285,-127</position>
<output>
<ID>OUT_0</ID>613 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>739</ID>
<type>GA_LED</type>
<position>300.5,-228</position>
<input>
<ID>N_in0</ID>614 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455,-138,455,-134</points>
<intersection>-138 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>455,-138,456,-138</points>
<connection>
<GID>490</GID>
<name>IN_1</name></connection>
<intersection>455 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>431.5,-134,455,-134</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>455 0</intersection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>460,-139,461,-139</points>
<connection>
<GID>490</GID>
<name>OUT</name></connection>
<connection>
<GID>462</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>455,-148,456,-148</points>
<connection>
<GID>485</GID>
<name>OUT</name></connection>
<connection>
<GID>463</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>447.5,-170.5,449.5,-170.5</points>
<connection>
<GID>465</GID>
<name>OUT</name></connection>
<connection>
<GID>464</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449.5,-186,449.5,-179.5</points>
<connection>
<GID>466</GID>
<name>IN_2</name></connection>
<intersection>-186 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-186,449.5,-186</points>
<connection>
<GID>469</GID>
<name>OUT</name></connection>
<intersection>449.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448.5,-181,448.5,-177.5</points>
<intersection>-181 2</intersection>
<intersection>-177.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>448.5,-177.5,449.5,-177.5</points>
<connection>
<GID>466</GID>
<name>IN_1</name></connection>
<intersection>448.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-181,448.5,-181</points>
<connection>
<GID>468</GID>
<name>OUT</name></connection>
<intersection>448.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>447.5,-175.5,449.5,-175.5</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<connection>
<GID>467</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>381,-90.5,382,-90.5</points>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<intersection>381 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>381,-91.5,381,-90.5</points>
<connection>
<GID>496</GID>
<name>OUT_0</name></connection>
<intersection>-90.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>455.5,-169.5,456.5,-169.5</points>
<connection>
<GID>470</GID>
<name>IN_0</name></connection>
<connection>
<GID>464</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432.5,-169.5,441.5,-169.5</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<intersection>439 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>439,-180,439,-169.5</points>
<intersection>-180 31</intersection>
<intersection>-174.5 29</intersection>
<intersection>-169.5 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>439,-174.5,441.5,-174.5</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<intersection>439 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>439,-180,441.5,-180</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>439 28</intersection></hsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436.5,-185,436.5,-171.5</points>
<intersection>-185 1</intersection>
<intersection>-176.5 4</intersection>
<intersection>-172.5 6</intersection>
<intersection>-171.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>436.5,-185,441.5,-185</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>436.5,-171.5,441.5,-171.5</points>
<connection>
<GID>465</GID>
<name>IN_1</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>436.5,-176.5,441.5,-176.5</points>
<connection>
<GID>467</GID>
<name>IN_1</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>432.5,-172.5,436.5,-172.5</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>441,-182,441.5,-182</points>
<connection>
<GID>471</GID>
<name>OUT_0</name></connection>
<connection>
<GID>468</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>441,-187,441.5,-187</points>
<connection>
<GID>472</GID>
<name>OUT_0</name></connection>
<connection>
<GID>469</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432,-166.5,449.5,-166.5</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>434.5 5</intersection>
<intersection>449.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>449.5,-168.5,449.5,-166.5</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<intersection>-166.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>434.5,-187,434.5,-166.5</points>
<intersection>-187 6</intersection>
<intersection>-182 8</intersection>
<intersection>-166.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>434.5,-187,437,-187</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<intersection>434.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>434.5,-182,437,-182</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<intersection>434.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458.5,-166,458.5,-160.5</points>
<connection>
<GID>470</GID>
<name>SEL_0</name></connection>
<intersection>-160.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432,-160.5,458.5,-160.5</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<intersection>458.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455.5,-167.5,455.5,-163.5</points>
<intersection>-167.5 1</intersection>
<intersection>-163.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>455.5,-167.5,456.5,-167.5</points>
<connection>
<GID>470</GID>
<name>IN_1</name></connection>
<intersection>455.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>432,-163.5,455.5,-163.5</points>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<intersection>455.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>460.5,-168.5,462,-168.5</points>
<connection>
<GID>470</GID>
<name>OUT</name></connection>
<connection>
<GID>478</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>455.5,-177.5,456.5,-177.5</points>
<connection>
<GID>466</GID>
<name>OUT</name></connection>
<connection>
<GID>479</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,-165.5,289,-163.5</points>
<intersection>-165.5 1</intersection>
<intersection>-163.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289,-165.5,290,-165.5</points>
<connection>
<GID>610</GID>
<name>IN_0</name></connection>
<intersection>289 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>287,-163.5,289,-163.5</points>
<connection>
<GID>613</GID>
<name>OUT_2</name></connection>
<intersection>289 0</intersection></hsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>446,-79.5,448,-79.5</points>
<connection>
<GID>499</GID>
<name>OUT</name></connection>
<connection>
<GID>498</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448,-95,448,-88.5</points>
<connection>
<GID>500</GID>
<name>IN_2</name></connection>
<intersection>-95 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>446,-95,448,-95</points>
<connection>
<GID>503</GID>
<name>OUT</name></connection>
<intersection>448 0</intersection></hsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>447,-90,447,-86.5</points>
<intersection>-90 2</intersection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>447,-86.5,448,-86.5</points>
<connection>
<GID>500</GID>
<name>IN_1</name></connection>
<intersection>447 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>446,-90,447,-90</points>
<connection>
<GID>502</GID>
<name>OUT</name></connection>
<intersection>447 0</intersection></hsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>446,-84.5,448,-84.5</points>
<connection>
<GID>500</GID>
<name>IN_0</name></connection>
<connection>
<GID>501</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>373,-79.5,375,-79.5</points>
<connection>
<GID>518</GID>
<name>IN_1</name></connection>
<connection>
<GID>519</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375,-95,375,-88.5</points>
<connection>
<GID>520</GID>
<name>IN_2</name></connection>
<intersection>-95 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>373,-95,375,-95</points>
<connection>
<GID>523</GID>
<name>OUT</name></connection>
<intersection>375 0</intersection></hsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374,-90,374,-86.5</points>
<intersection>-90 2</intersection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>374,-86.5,375,-86.5</points>
<connection>
<GID>520</GID>
<name>IN_1</name></connection>
<intersection>374 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>373,-90,374,-90</points>
<connection>
<GID>522</GID>
<name>OUT</name></connection>
<intersection>374 0</intersection></hsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>373,-84.5,375,-84.5</points>
<connection>
<GID>520</GID>
<name>IN_0</name></connection>
<connection>
<GID>521</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>381,-78.5,382,-78.5</points>
<connection>
<GID>518</GID>
<name>OUT</name></connection>
<connection>
<GID>524</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>454,-78.5,455,-78.5</points>
<connection>
<GID>504</GID>
<name>IN_0</name></connection>
<connection>
<GID>498</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>431,-78.5,440,-78.5</points>
<connection>
<GID>499</GID>
<name>IN_0</name></connection>
<connection>
<GID>510</GID>
<name>IN_0</name></connection>
<intersection>437.5 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>437.5,-89,437.5,-78.5</points>
<intersection>-89 31</intersection>
<intersection>-83.5 29</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>437.5,-83.5,440,-83.5</points>
<connection>
<GID>501</GID>
<name>IN_0</name></connection>
<intersection>437.5 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>437.5,-89,440,-89</points>
<connection>
<GID>502</GID>
<name>IN_0</name></connection>
<intersection>437.5 28</intersection></hsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>358,-78.5,367,-78.5</points>
<connection>
<GID>519</GID>
<name>IN_0</name></connection>
<connection>
<GID>557</GID>
<name>IN_0</name></connection>
<intersection>364.5 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>364.5,-89,364.5,-78.5</points>
<intersection>-89 31</intersection>
<intersection>-83.5 29</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>364.5,-83.5,367,-83.5</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<intersection>364.5 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>364.5,-89,367,-89</points>
<connection>
<GID>522</GID>
<name>IN_0</name></connection>
<intersection>364.5 28</intersection></hsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>435,-94,435,-80.5</points>
<intersection>-94 1</intersection>
<intersection>-85.5 4</intersection>
<intersection>-81.5 6</intersection>
<intersection>-80.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>435,-94,440,-94</points>
<connection>
<GID>503</GID>
<name>IN_0</name></connection>
<intersection>435 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>435,-80.5,440,-80.5</points>
<connection>
<GID>499</GID>
<name>IN_1</name></connection>
<intersection>435 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>435,-85.5,440,-85.5</points>
<connection>
<GID>501</GID>
<name>IN_1</name></connection>
<intersection>435 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>431,-81.5,435,-81.5</points>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<intersection>435 0</intersection></hsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>362,-94,362,-80.5</points>
<intersection>-94 1</intersection>
<intersection>-85.5 4</intersection>
<intersection>-81.5 6</intersection>
<intersection>-80.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>362,-94,367,-94</points>
<connection>
<GID>523</GID>
<name>IN_0</name></connection>
<intersection>362 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>362,-80.5,367,-80.5</points>
<connection>
<GID>519</GID>
<name>IN_1</name></connection>
<intersection>362 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>362,-85.5,367,-85.5</points>
<connection>
<GID>521</GID>
<name>IN_1</name></connection>
<intersection>362 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>358,-81.5,362,-81.5</points>
<connection>
<GID>558</GID>
<name>IN_0</name></connection>
<intersection>362 0</intersection></hsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>366.5,-91,367,-91</points>
<connection>
<GID>522</GID>
<name>IN_1</name></connection>
<connection>
<GID>530</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>366.5,-96,367,-96</points>
<connection>
<GID>523</GID>
<name>IN_1</name></connection>
<connection>
<GID>531</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>439.5,-91,440,-91</points>
<connection>
<GID>505</GID>
<name>OUT_0</name></connection>
<connection>
<GID>502</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>439.5,-96,440,-96</points>
<connection>
<GID>506</GID>
<name>OUT_0</name></connection>
<connection>
<GID>503</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>430.5,-75.5,448,-75.5</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>433 5</intersection>
<intersection>448 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>448,-77.5,448,-75.5</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>433,-96,433,-75.5</points>
<intersection>-96 6</intersection>
<intersection>-91 8</intersection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>433,-96,435.5,-96</points>
<connection>
<GID>506</GID>
<name>IN_0</name></connection>
<intersection>433 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>433,-91,435.5,-91</points>
<connection>
<GID>505</GID>
<name>IN_0</name></connection>
<intersection>433 5</intersection></hsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457,-75,457,-69.5</points>
<connection>
<GID>504</GID>
<name>SEL_0</name></connection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>430.5,-69.5,457,-69.5</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<intersection>457 0</intersection></hsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454,-76.5,454,-72.5</points>
<intersection>-76.5 1</intersection>
<intersection>-72.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>454,-76.5,455,-76.5</points>
<connection>
<GID>504</GID>
<name>IN_1</name></connection>
<intersection>454 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>430.5,-72.5,454,-72.5</points>
<connection>
<GID>508</GID>
<name>IN_0</name></connection>
<intersection>454 0</intersection></hsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>357.5,-75.5,375,-75.5</points>
<connection>
<GID>556</GID>
<name>IN_0</name></connection>
<intersection>360 5</intersection>
<intersection>375 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>375,-77.5,375,-75.5</points>
<connection>
<GID>518</GID>
<name>IN_0</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>360,-96,360,-75.5</points>
<intersection>-96 6</intersection>
<intersection>-91 8</intersection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>360,-96,362.5,-96</points>
<connection>
<GID>531</GID>
<name>IN_0</name></connection>
<intersection>360 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>360,-91,362.5,-91</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<intersection>360 5</intersection></hsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>459,-77.5,460,-77.5</points>
<connection>
<GID>504</GID>
<name>OUT</name></connection>
<connection>
<GID>512</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384,-75,384,-69.5</points>
<connection>
<GID>524</GID>
<name>SEL_0</name></connection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>357.5,-69.5,384,-69.5</points>
<connection>
<GID>553</GID>
<name>IN_0</name></connection>
<intersection>384 0</intersection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>381,-76.5,381,-72.5</points>
<intersection>-76.5 1</intersection>
<intersection>-72.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381,-76.5,382,-76.5</points>
<connection>
<GID>524</GID>
<name>IN_1</name></connection>
<intersection>381 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357.5,-72.5,381,-72.5</points>
<connection>
<GID>555</GID>
<name>IN_0</name></connection>
<intersection>381 0</intersection></hsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>386,-77.5,387,-77.5</points>
<connection>
<GID>524</GID>
<name>OUT</name></connection>
<connection>
<GID>559</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>381,-86.5,382,-86.5</points>
<connection>
<GID>520</GID>
<name>OUT</name></connection>
<connection>
<GID>560</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>454,-86.5,455,-86.5</points>
<connection>
<GID>500</GID>
<name>OUT</name></connection>
<connection>
<GID>513</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>373.5,-109,375.5,-109</points>
<connection>
<GID>564</GID>
<name>OUT</name></connection>
<connection>
<GID>563</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375.5,-124.5,375.5,-118</points>
<connection>
<GID>565</GID>
<name>IN_2</name></connection>
<intersection>-124.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>373.5,-124.5,375.5,-124.5</points>
<connection>
<GID>568</GID>
<name>OUT</name></connection>
<intersection>375.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374.5,-119.5,374.5,-116</points>
<intersection>-119.5 2</intersection>
<intersection>-116 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>374.5,-116,375.5,-116</points>
<connection>
<GID>565</GID>
<name>IN_1</name></connection>
<intersection>374.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>373.5,-119.5,374.5,-119.5</points>
<connection>
<GID>567</GID>
<name>OUT</name></connection>
<intersection>374.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>373.5,-114,375.5,-114</points>
<connection>
<GID>565</GID>
<name>IN_0</name></connection>
<connection>
<GID>566</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>381.5,-108,382.5,-108</points>
<connection>
<GID>569</GID>
<name>IN_0</name></connection>
<connection>
<GID>563</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>358.5,-108,367.5,-108</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<connection>
<GID>575</GID>
<name>IN_0</name></connection>
<intersection>365 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>365,-118.5,365,-108</points>
<intersection>-118.5 31</intersection>
<intersection>-113 29</intersection>
<intersection>-108 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>365,-113,367.5,-113</points>
<connection>
<GID>566</GID>
<name>IN_0</name></connection>
<intersection>365 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>365,-118.5,367.5,-118.5</points>
<connection>
<GID>567</GID>
<name>IN_0</name></connection>
<intersection>365 28</intersection></hsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>362.5,-123.5,362.5,-110</points>
<intersection>-123.5 1</intersection>
<intersection>-115 4</intersection>
<intersection>-111 6</intersection>
<intersection>-110 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>362.5,-123.5,367.5,-123.5</points>
<connection>
<GID>568</GID>
<name>IN_0</name></connection>
<intersection>362.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>362.5,-110,367.5,-110</points>
<connection>
<GID>564</GID>
<name>IN_1</name></connection>
<intersection>362.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>362.5,-115,367.5,-115</points>
<connection>
<GID>566</GID>
<name>IN_1</name></connection>
<intersection>362.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>358.5,-111,362.5,-111</points>
<connection>
<GID>576</GID>
<name>IN_0</name></connection>
<intersection>362.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>367,-120.5,367.5,-120.5</points>
<connection>
<GID>570</GID>
<name>OUT_0</name></connection>
<connection>
<GID>567</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>367,-125.5,367.5,-125.5</points>
<connection>
<GID>571</GID>
<name>OUT_0</name></connection>
<connection>
<GID>568</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>358,-105,375.5,-105</points>
<connection>
<GID>574</GID>
<name>IN_0</name></connection>
<intersection>360.5 5</intersection>
<intersection>375.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>375.5,-107,375.5,-105</points>
<connection>
<GID>563</GID>
<name>IN_0</name></connection>
<intersection>-105 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>360.5,-125.5,360.5,-105</points>
<intersection>-125.5 6</intersection>
<intersection>-120.5 8</intersection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>360.5,-125.5,363,-125.5</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>360.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>360.5,-120.5,363,-120.5</points>
<connection>
<GID>570</GID>
<name>IN_0</name></connection>
<intersection>360.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384.5,-104.5,384.5,-99</points>
<connection>
<GID>569</GID>
<name>SEL_0</name></connection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>358,-99,384.5,-99</points>
<connection>
<GID>572</GID>
<name>IN_0</name></connection>
<intersection>384.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>381.5,-106,381.5,-102</points>
<intersection>-106 1</intersection>
<intersection>-102 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381.5,-106,382.5,-106</points>
<connection>
<GID>569</GID>
<name>IN_1</name></connection>
<intersection>381.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>358,-102,381.5,-102</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<intersection>381.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>386.5,-107,388,-107</points>
<connection>
<GID>569</GID>
<name>OUT</name></connection>
<connection>
<GID>577</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>381.5,-116,382.5,-116</points>
<connection>
<GID>565</GID>
<name>OUT</name></connection>
<connection>
<GID>578</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>446.5,-109,448.5,-109</points>
<connection>
<GID>515</GID>
<name>OUT</name></connection>
<connection>
<GID>514</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448.5,-124.5,448.5,-118</points>
<connection>
<GID>517</GID>
<name>IN_2</name></connection>
<intersection>-124.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>446.5,-124.5,448.5,-124.5</points>
<connection>
<GID>527</GID>
<name>OUT</name></connection>
<intersection>448.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>447.5,-119.5,447.5,-116</points>
<intersection>-119.5 2</intersection>
<intersection>-116 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>447.5,-116,448.5,-116</points>
<connection>
<GID>517</GID>
<name>IN_1</name></connection>
<intersection>447.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>446.5,-119.5,447.5,-119.5</points>
<connection>
<GID>526</GID>
<name>OUT</name></connection>
<intersection>447.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>446.5,-114,448.5,-114</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<connection>
<GID>525</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>454.5,-108,455.5,-108</points>
<connection>
<GID>528</GID>
<name>IN_0</name></connection>
<connection>
<GID>514</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>431.5,-108,440.5,-108</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<connection>
<GID>536</GID>
<name>IN_0</name></connection>
<intersection>438 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>438,-118.5,438,-108</points>
<intersection>-118.5 31</intersection>
<intersection>-113 29</intersection>
<intersection>-108 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>438,-113,440.5,-113</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<intersection>438 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>438,-118.5,440.5,-118.5</points>
<connection>
<GID>526</GID>
<name>IN_0</name></connection>
<intersection>438 28</intersection></hsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>435.5,-123.5,435.5,-110</points>
<intersection>-123.5 1</intersection>
<intersection>-115 4</intersection>
<intersection>-111 6</intersection>
<intersection>-110 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>435.5,-123.5,440.5,-123.5</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<intersection>435.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>435.5,-110,440.5,-110</points>
<connection>
<GID>515</GID>
<name>IN_1</name></connection>
<intersection>435.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>435.5,-115,440.5,-115</points>
<connection>
<GID>525</GID>
<name>IN_1</name></connection>
<intersection>435.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>431.5,-111,435.5,-111</points>
<connection>
<GID>537</GID>
<name>IN_0</name></connection>
<intersection>435.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440,-120.5,440.5,-120.5</points>
<connection>
<GID>529</GID>
<name>OUT_0</name></connection>
<connection>
<GID>526</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440,-125.5,440.5,-125.5</points>
<connection>
<GID>532</GID>
<name>OUT_0</name></connection>
<connection>
<GID>527</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>431,-105,448.5,-105</points>
<connection>
<GID>535</GID>
<name>IN_0</name></connection>
<intersection>433.5 5</intersection>
<intersection>448.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>448.5,-107,448.5,-105</points>
<connection>
<GID>514</GID>
<name>IN_0</name></connection>
<intersection>-105 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>433.5,-125.5,433.5,-105</points>
<intersection>-125.5 6</intersection>
<intersection>-120.5 8</intersection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>433.5,-125.5,436,-125.5</points>
<connection>
<GID>532</GID>
<name>IN_0</name></connection>
<intersection>433.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>433.5,-120.5,436,-120.5</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<intersection>433.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457.5,-104.5,457.5,-99</points>
<connection>
<GID>528</GID>
<name>SEL_0</name></connection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>431,-99,457.5,-99</points>
<connection>
<GID>533</GID>
<name>IN_0</name></connection>
<intersection>457.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454.5,-106,454.5,-102</points>
<intersection>-106 1</intersection>
<intersection>-102 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>454.5,-106,455.5,-106</points>
<connection>
<GID>528</GID>
<name>IN_1</name></connection>
<intersection>454.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>431,-102,454.5,-102</points>
<connection>
<GID>534</GID>
<name>IN_0</name></connection>
<intersection>454.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>459.5,-107,461,-107</points>
<connection>
<GID>528</GID>
<name>OUT</name></connection>
<connection>
<GID>538</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>454.5,-116,455.5,-116</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<connection>
<GID>517</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,-168.5,288.5,-164.5</points>
<intersection>-168.5 1</intersection>
<intersection>-164.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288.5,-168.5,290,-168.5</points>
<connection>
<GID>611</GID>
<name>IN_0</name></connection>
<intersection>288.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>287,-164.5,288.5,-164.5</points>
<connection>
<GID>613</GID>
<name>OUT_3</name></connection>
<intersection>288.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>375.5,-267.5,377.5,-267.5</points>
<connection>
<GID>629</GID>
<name>OUT</name></connection>
<connection>
<GID>626</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>466</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>377.5,-283,377.5,-276.5</points>
<connection>
<GID>630</GID>
<name>IN_2</name></connection>
<intersection>-283 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>375.5,-283,377.5,-283</points>
<connection>
<GID>645</GID>
<name>OUT</name></connection>
<intersection>377.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>376.5,-278,376.5,-274.5</points>
<intersection>-278 2</intersection>
<intersection>-274.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>376.5,-274.5,377.5,-274.5</points>
<connection>
<GID>630</GID>
<name>IN_1</name></connection>
<intersection>376.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375.5,-278,376.5,-278</points>
<connection>
<GID>643</GID>
<name>OUT</name></connection>
<intersection>376.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>375,-272.5,377.5,-272.5</points>
<connection>
<GID>630</GID>
<name>IN_0</name></connection>
<connection>
<GID>638</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>469</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>383.5,-266.5,384.5,-266.5</points>
<connection>
<GID>626</GID>
<name>OUT</name></connection>
<connection>
<GID>647</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>360.5,-266.5,369.5,-266.5</points>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<connection>
<GID>540</GID>
<name>IN_0</name></connection>
<intersection>367 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>367,-277,367,-266.5</points>
<intersection>-277 31</intersection>
<intersection>-271.5 29</intersection>
<intersection>-266.5 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>367,-271.5,369,-271.5</points>
<connection>
<GID>638</GID>
<name>IN_0</name></connection>
<intersection>367 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>367,-277,369.5,-277</points>
<connection>
<GID>643</GID>
<name>IN_0</name></connection>
<intersection>367 28</intersection></hsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>364.5,-282,364.5,-268.5</points>
<intersection>-282 1</intersection>
<intersection>-273.5 4</intersection>
<intersection>-269.5 6</intersection>
<intersection>-268.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>364.5,-282,369.5,-282</points>
<connection>
<GID>645</GID>
<name>IN_0</name></connection>
<intersection>364.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>364.5,-268.5,369.5,-268.5</points>
<connection>
<GID>629</GID>
<name>IN_1</name></connection>
<intersection>364.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>364.5,-273.5,369,-273.5</points>
<connection>
<GID>638</GID>
<name>IN_1</name></connection>
<intersection>364.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>360.5,-269.5,364.5,-269.5</points>
<connection>
<GID>541</GID>
<name>IN_0</name></connection>
<intersection>364.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>369,-279,369.5,-279</points>
<connection>
<GID>649</GID>
<name>OUT_0</name></connection>
<connection>
<GID>643</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>369,-284,369.5,-284</points>
<connection>
<GID>652</GID>
<name>OUT_0</name></connection>
<connection>
<GID>645</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>360,-263.5,377.5,-263.5</points>
<connection>
<GID>660</GID>
<name>IN_0</name></connection>
<intersection>362.5 5</intersection>
<intersection>377.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>377.5,-265.5,377.5,-263.5</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>-263.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>362.5,-284,362.5,-263.5</points>
<intersection>-284 6</intersection>
<intersection>-279 8</intersection>
<intersection>-263.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>362.5,-284,365,-284</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<intersection>362.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>362.5,-279,365,-279</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<intersection>362.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>386.5,-263,386.5,-257.5</points>
<connection>
<GID>647</GID>
<name>SEL_0</name></connection>
<intersection>-257.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360,-257.5,386.5,-257.5</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<intersection>386.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>383.5,-264.5,383.5,-260.5</points>
<intersection>-264.5 1</intersection>
<intersection>-260.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>383.5,-264.5,384.5,-264.5</points>
<connection>
<GID>647</GID>
<name>IN_1</name></connection>
<intersection>383.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>360,-260.5,383.5,-260.5</points>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<intersection>383.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>388.5,-265.5,389.5,-265.5</points>
<connection>
<GID>647</GID>
<name>OUT</name></connection>
<connection>
<GID>542</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>383.5,-274.5,384.5,-274.5</points>
<connection>
<GID>630</GID>
<name>OUT</name></connection>
<connection>
<GID>543</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>376,-297,378,-297</points>
<connection>
<GID>545</GID>
<name>OUT</name></connection>
<connection>
<GID>544</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>378,-312.5,378,-306</points>
<connection>
<GID>546</GID>
<name>IN_2</name></connection>
<intersection>-312.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>376,-312.5,378,-312.5</points>
<connection>
<GID>549</GID>
<name>OUT</name></connection>
<intersection>378 0</intersection></hsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>377,-307.5,377,-304</points>
<intersection>-307.5 2</intersection>
<intersection>-304 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>377,-304,378,-304</points>
<connection>
<GID>546</GID>
<name>IN_1</name></connection>
<intersection>377 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>376,-307.5,377,-307.5</points>
<connection>
<GID>548</GID>
<name>OUT</name></connection>
<intersection>377 0</intersection></hsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>14</ID>
<points>376,-302.5,376,-302</points>
<connection>
<GID>547</GID>
<name>OUT</name></connection>
<intersection>-302 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>376,-302,378,-302</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<intersection>376 14</intersection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>384,-296,385,-296</points>
<connection>
<GID>544</GID>
<name>OUT</name></connection>
<connection>
<GID>550</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>361,-296,370,-296</points>
<connection>
<GID>545</GID>
<name>IN_0</name></connection>
<connection>
<GID>579</GID>
<name>IN_0</name></connection>
<intersection>361 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>361,-306.5,361,-296</points>
<intersection>-306.5 31</intersection>
<intersection>-301.5 29</intersection>
<intersection>-296 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>361,-301.5,370,-301.5</points>
<connection>
<GID>547</GID>
<name>IN_0</name></connection>
<intersection>361 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>361,-306.5,370,-306.5</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<intersection>361 28</intersection></hsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>365,-311.5,365,-298</points>
<intersection>-311.5 1</intersection>
<intersection>-303.5 4</intersection>
<intersection>-299 6</intersection>
<intersection>-298 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>365,-311.5,370,-311.5</points>
<connection>
<GID>549</GID>
<name>IN_0</name></connection>
<intersection>365 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>365,-298,370,-298</points>
<connection>
<GID>545</GID>
<name>IN_1</name></connection>
<intersection>365 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>365,-303.5,370,-303.5</points>
<connection>
<GID>547</GID>
<name>IN_1</name></connection>
<intersection>365 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>361,-299,365,-299</points>
<connection>
<GID>581</GID>
<name>IN_0</name></connection>
<intersection>365 0</intersection></hsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>369.5,-308.5,370,-308.5</points>
<connection>
<GID>551</GID>
<name>OUT_0</name></connection>
<connection>
<GID>548</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>369.5,-313.5,370,-313.5</points>
<connection>
<GID>552</GID>
<name>OUT_0</name></connection>
<connection>
<GID>549</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>360.5,-293,378,-293</points>
<connection>
<GID>562</GID>
<name>IN_0</name></connection>
<intersection>363 5</intersection>
<intersection>378 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>378,-295,378,-293</points>
<connection>
<GID>544</GID>
<name>IN_0</name></connection>
<intersection>-293 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>363,-313.5,363,-293</points>
<intersection>-313.5 6</intersection>
<intersection>-308.5 8</intersection>
<intersection>-293 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>363,-313.5,365.5,-313.5</points>
<connection>
<GID>552</GID>
<name>IN_0</name></connection>
<intersection>363 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>363,-308.5,365.5,-308.5</points>
<connection>
<GID>551</GID>
<name>IN_0</name></connection>
<intersection>363 5</intersection></hsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>387,-292.5,387,-287</points>
<connection>
<GID>550</GID>
<name>SEL_0</name></connection>
<intersection>-287 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360.5,-287,387,-287</points>
<connection>
<GID>554</GID>
<name>IN_0</name></connection>
<intersection>387 0</intersection></hsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384,-294,384,-290</points>
<intersection>-294 1</intersection>
<intersection>-290 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384,-294,385,-294</points>
<connection>
<GID>550</GID>
<name>IN_1</name></connection>
<intersection>384 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>360.5,-290,384,-290</points>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<intersection>384 0</intersection></hsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>389,-295,390.5,-295</points>
<connection>
<GID>550</GID>
<name>OUT</name></connection>
<connection>
<GID>583</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>384,-304,385,-304</points>
<connection>
<GID>546</GID>
<name>OUT</name></connection>
<connection>
<GID>585</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,-161.5,289,-159.5</points>
<intersection>-161.5 1</intersection>
<intersection>-159.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287,-161.5,289,-161.5</points>
<connection>
<GID>613</GID>
<name>OUT_0</name></connection>
<intersection>289 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>289,-159.5,290,-159.5</points>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<intersection>289 0</intersection></hsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>448.5,-267.5,450.5,-267.5</points>
<connection>
<GID>614</GID>
<name>OUT</name></connection>
<connection>
<GID>612</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>450.5,-283,450.5,-276.5</points>
<connection>
<GID>615</GID>
<name>IN_2</name></connection>
<intersection>-283 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>448.5,-283,450.5,-283</points>
<connection>
<GID>619</GID>
<name>OUT</name></connection>
<intersection>450.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449.5,-278,449.5,-274.5</points>
<intersection>-278 2</intersection>
<intersection>-274.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>449.5,-274.5,450.5,-274.5</points>
<connection>
<GID>615</GID>
<name>IN_1</name></connection>
<intersection>449.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448.5,-278,449.5,-278</points>
<connection>
<GID>618</GID>
<name>OUT</name></connection>
<intersection>449.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>448.5,-272.5,450.5,-272.5</points>
<connection>
<GID>615</GID>
<name>IN_0</name></connection>
<connection>
<GID>617</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>456.5,-266.5,457.5,-266.5</points>
<connection>
<GID>612</GID>
<name>OUT</name></connection>
<connection>
<GID>620</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>433.5,-266.5,442.5,-266.5</points>
<connection>
<GID>614</GID>
<name>IN_0</name></connection>
<connection>
<GID>587</GID>
<name>IN_0</name></connection>
<intersection>440 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>440,-277,440,-266.5</points>
<intersection>-277 31</intersection>
<intersection>-271.5 29</intersection>
<intersection>-266.5 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>440,-271.5,442.5,-271.5</points>
<connection>
<GID>617</GID>
<name>IN_0</name></connection>
<intersection>440 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>440,-277,442.5,-277</points>
<connection>
<GID>618</GID>
<name>IN_0</name></connection>
<intersection>440 28</intersection></hsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>437.5,-282,437.5,-268.5</points>
<intersection>-282 1</intersection>
<intersection>-273.5 4</intersection>
<intersection>-269.5 6</intersection>
<intersection>-268.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>437.5,-282,442.5,-282</points>
<connection>
<GID>619</GID>
<name>IN_0</name></connection>
<intersection>437.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>437.5,-268.5,442.5,-268.5</points>
<connection>
<GID>614</GID>
<name>IN_1</name></connection>
<intersection>437.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>437.5,-273.5,442.5,-273.5</points>
<connection>
<GID>617</GID>
<name>IN_1</name></connection>
<intersection>437.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>433.5,-269.5,437.5,-269.5</points>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<intersection>437.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>442,-279,442.5,-279</points>
<connection>
<GID>621</GID>
<name>OUT_0</name></connection>
<connection>
<GID>618</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>442,-284,442.5,-284</points>
<connection>
<GID>622</GID>
<name>OUT_0</name></connection>
<connection>
<GID>619</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>433,-263.5,450.5,-263.5</points>
<connection>
<GID>632</GID>
<name>IN_0</name></connection>
<intersection>435.5 5</intersection>
<intersection>450.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>450.5,-265.5,450.5,-263.5</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<intersection>-263.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>435.5,-284,435.5,-263.5</points>
<intersection>-284 6</intersection>
<intersection>-279 8</intersection>
<intersection>-263.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>435.5,-284,438,-284</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<intersection>435.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>435.5,-279,438,-279</points>
<connection>
<GID>621</GID>
<name>IN_0</name></connection>
<intersection>435.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459.5,-263,459.5,-257.5</points>
<connection>
<GID>620</GID>
<name>SEL_0</name></connection>
<intersection>-257.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>433,-257.5,459.5,-257.5</points>
<connection>
<GID>624</GID>
<name>IN_0</name></connection>
<intersection>459.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456.5,-264.5,456.5,-260.5</points>
<intersection>-264.5 1</intersection>
<intersection>-260.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>456.5,-264.5,457.5,-264.5</points>
<connection>
<GID>620</GID>
<name>IN_1</name></connection>
<intersection>456.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>433,-260.5,456.5,-260.5</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<intersection>456.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>461.5,-265.5,462.5,-265.5</points>
<connection>
<GID>620</GID>
<name>OUT</name></connection>
<connection>
<GID>591</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>456.5,-274.5,457.5,-274.5</points>
<connection>
<GID>615</GID>
<name>OUT</name></connection>
<connection>
<GID>593</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>449,-297,451,-297</points>
<connection>
<GID>595</GID>
<name>OUT</name></connection>
<connection>
<GID>594</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>451,-312.5,451,-306</points>
<connection>
<GID>596</GID>
<name>IN_2</name></connection>
<intersection>-312.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>449,-312.5,451,-312.5</points>
<connection>
<GID>599</GID>
<name>OUT</name></connection>
<intersection>451 0</intersection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>450,-307.5,450,-304</points>
<intersection>-307.5 2</intersection>
<intersection>-304 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>450,-304,451,-304</points>
<connection>
<GID>596</GID>
<name>IN_1</name></connection>
<intersection>450 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>449,-307.5,450,-307.5</points>
<connection>
<GID>598</GID>
<name>OUT</name></connection>
<intersection>450 0</intersection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<vsegment>
<ID>14</ID>
<points>449,-302.5,449,-302</points>
<connection>
<GID>597</GID>
<name>OUT</name></connection>
<intersection>-302 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>449,-302,451,-302</points>
<connection>
<GID>596</GID>
<name>IN_0</name></connection>
<intersection>449 14</intersection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>274,-161,279,-161</points>
<connection>
<GID>613</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>616</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>457,-296,458,-296</points>
<connection>
<GID>594</GID>
<name>OUT</name></connection>
<connection>
<GID>600</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>434,-296,443,-296</points>
<connection>
<GID>595</GID>
<name>IN_0</name></connection>
<connection>
<GID>606</GID>
<name>IN_0</name></connection>
<intersection>434 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>434,-306.5,434,-296</points>
<intersection>-306.5 31</intersection>
<intersection>-301.5 29</intersection>
<intersection>-296 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>434,-301.5,443,-301.5</points>
<connection>
<GID>597</GID>
<name>IN_0</name></connection>
<intersection>434 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>434,-306.5,443,-306.5</points>
<connection>
<GID>598</GID>
<name>IN_0</name></connection>
<intersection>434 28</intersection></hsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>438,-311.5,438,-298</points>
<intersection>-311.5 1</intersection>
<intersection>-303.5 4</intersection>
<intersection>-299 6</intersection>
<intersection>-298 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>438,-311.5,443,-311.5</points>
<connection>
<GID>599</GID>
<name>IN_0</name></connection>
<intersection>438 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>438,-298,443,-298</points>
<connection>
<GID>595</GID>
<name>IN_1</name></connection>
<intersection>438 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>438,-303.5,443,-303.5</points>
<connection>
<GID>597</GID>
<name>IN_1</name></connection>
<intersection>438 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>434,-299,438,-299</points>
<connection>
<GID>607</GID>
<name>IN_0</name></connection>
<intersection>438 0</intersection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>442.5,-308.5,443,-308.5</points>
<connection>
<GID>601</GID>
<name>OUT_0</name></connection>
<connection>
<GID>598</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>442.5,-313.5,443,-313.5</points>
<connection>
<GID>602</GID>
<name>OUT_0</name></connection>
<connection>
<GID>599</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>433.5,-293,451,-293</points>
<connection>
<GID>605</GID>
<name>IN_0</name></connection>
<intersection>436 5</intersection>
<intersection>451 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>451,-295,451,-293</points>
<connection>
<GID>594</GID>
<name>IN_0</name></connection>
<intersection>-293 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>436,-313.5,436,-293</points>
<intersection>-313.5 6</intersection>
<intersection>-308.5 8</intersection>
<intersection>-293 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>436,-313.5,438.5,-313.5</points>
<connection>
<GID>602</GID>
<name>IN_0</name></connection>
<intersection>436 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>436,-308.5,438.5,-308.5</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<intersection>436 5</intersection></hsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>460,-292.5,460,-287</points>
<connection>
<GID>600</GID>
<name>SEL_0</name></connection>
<intersection>-287 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>433.5,-287,460,-287</points>
<connection>
<GID>603</GID>
<name>IN_0</name></connection>
<intersection>460 0</intersection></hsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457,-294,457,-290</points>
<intersection>-294 1</intersection>
<intersection>-290 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>457,-294,458,-294</points>
<connection>
<GID>600</GID>
<name>IN_1</name></connection>
<intersection>457 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>433.5,-290,457,-290</points>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<intersection>457 0</intersection></hsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>462,-295,463.5,-295</points>
<connection>
<GID>600</GID>
<name>OUT</name></connection>
<connection>
<GID>608</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-160,276,-157.5</points>
<intersection>-160 2</intersection>
<intersection>-157.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274,-157.5,276,-157.5</points>
<connection>
<GID>706</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-160,279,-160</points>
<connection>
<GID>613</GID>
<name>IN_B_2</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277,-159,277,-154.5</points>
<intersection>-159 2</intersection>
<intersection>-154.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274,-154.5,277,-154.5</points>
<connection>
<GID>708</GID>
<name>IN_0</name></connection>
<intersection>277 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277,-159,279,-159</points>
<connection>
<GID>613</GID>
<name>IN_B_1</name></connection>
<intersection>277 0</intersection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>447.5,-206,449.5,-206</points>
<connection>
<GID>634</GID>
<name>OUT</name></connection>
<connection>
<GID>633</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449.5,-221.5,449.5,-215</points>
<connection>
<GID>635</GID>
<name>IN_2</name></connection>
<intersection>-221.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-221.5,449.5,-221.5</points>
<connection>
<GID>639</GID>
<name>OUT</name></connection>
<intersection>449.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448.5,-216.5,448.5,-213</points>
<intersection>-216.5 2</intersection>
<intersection>-213 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>448.5,-213,449.5,-213</points>
<connection>
<GID>635</GID>
<name>IN_1</name></connection>
<intersection>448.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-216.5,448.5,-216.5</points>
<connection>
<GID>637</GID>
<name>OUT</name></connection>
<intersection>448.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>447.5,-211,449.5,-211</points>
<connection>
<GID>635</GID>
<name>IN_0</name></connection>
<connection>
<GID>636</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>374.5,-206,376.5,-206</points>
<connection>
<GID>662</GID>
<name>OUT</name></connection>
<connection>
<GID>661</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>376.5,-221.5,376.5,-215</points>
<connection>
<GID>663</GID>
<name>IN_2</name></connection>
<intersection>-221.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>374.5,-221.5,376.5,-221.5</points>
<connection>
<GID>666</GID>
<name>OUT</name></connection>
<intersection>376.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375.5,-216.5,375.5,-213</points>
<intersection>-216.5 2</intersection>
<intersection>-213 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375.5,-213,376.5,-213</points>
<connection>
<GID>663</GID>
<name>IN_1</name></connection>
<intersection>375.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>374.5,-216.5,375.5,-216.5</points>
<connection>
<GID>665</GID>
<name>OUT</name></connection>
<intersection>375.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>374.5,-211,376.5,-211</points>
<connection>
<GID>663</GID>
<name>IN_0</name></connection>
<connection>
<GID>664</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382.5,-205,383.5,-205</points>
<connection>
<GID>661</GID>
<name>OUT</name></connection>
<connection>
<GID>667</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>455.5,-205,456.5,-205</points>
<connection>
<GID>633</GID>
<name>OUT</name></connection>
<connection>
<GID>640</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432.5,-205,441.5,-205</points>
<connection>
<GID>634</GID>
<name>IN_0</name></connection>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<intersection>432.5 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>432.5,-215.5,432.5,-205</points>
<intersection>-215.5 31</intersection>
<intersection>-210 29</intersection>
<intersection>-205 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>432.5,-210,441.5,-210</points>
<connection>
<GID>636</GID>
<name>IN_0</name></connection>
<intersection>432.5 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>432.5,-215.5,441.5,-215.5</points>
<connection>
<GID>637</GID>
<name>IN_0</name></connection>
<intersection>432.5 28</intersection></hsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>359.5,-205,368.5,-205</points>
<connection>
<GID>662</GID>
<name>IN_0</name></connection>
<connection>
<GID>686</GID>
<name>IN_0</name></connection>
<intersection>359.5 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>359.5,-215.5,359.5,-205</points>
<intersection>-215.5 31</intersection>
<intersection>-210 29</intersection>
<intersection>-205 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>359.5,-210,368.5,-210</points>
<connection>
<GID>664</GID>
<name>IN_0</name></connection>
<intersection>359.5 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>359.5,-215.5,368.5,-215.5</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<intersection>359.5 28</intersection></hsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436.5,-220.5,436.5,-207</points>
<intersection>-220.5 1</intersection>
<intersection>-212 4</intersection>
<intersection>-208 6</intersection>
<intersection>-207 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>436.5,-220.5,441.5,-220.5</points>
<connection>
<GID>639</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>436.5,-207,441.5,-207</points>
<connection>
<GID>634</GID>
<name>IN_1</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>436.5,-212,441.5,-212</points>
<connection>
<GID>636</GID>
<name>IN_1</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>432.5,-208,436.5,-208</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363.5,-220.5,363.5,-207</points>
<intersection>-220.5 1</intersection>
<intersection>-212 4</intersection>
<intersection>-208 6</intersection>
<intersection>-207 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>363.5,-220.5,368.5,-220.5</points>
<connection>
<GID>666</GID>
<name>IN_0</name></connection>
<intersection>363.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>363.5,-207,368.5,-207</points>
<connection>
<GID>662</GID>
<name>IN_1</name></connection>
<intersection>363.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>363.5,-212,368.5,-212</points>
<connection>
<GID>664</GID>
<name>IN_1</name></connection>
<intersection>363.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>359.5,-208,363.5,-208</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<intersection>363.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>538</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>368,-217.5,368.5,-217.5</points>
<connection>
<GID>673</GID>
<name>OUT_0</name></connection>
<connection>
<GID>665</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>368,-222.5,368.5,-222.5</points>
<connection>
<GID>674</GID>
<name>OUT_0</name></connection>
<connection>
<GID>666</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>441,-217.5,441.5,-217.5</points>
<connection>
<GID>641</GID>
<name>OUT_0</name></connection>
<connection>
<GID>637</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>441,-222.5,441.5,-222.5</points>
<connection>
<GID>642</GID>
<name>OUT_0</name></connection>
<connection>
<GID>639</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432,-202,449.5,-202</points>
<connection>
<GID>648</GID>
<name>IN_0</name></connection>
<intersection>434.5 5</intersection>
<intersection>449.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>449.5,-204,449.5,-202</points>
<connection>
<GID>633</GID>
<name>IN_0</name></connection>
<intersection>-202 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>434.5,-222.5,434.5,-202</points>
<intersection>-222.5 6</intersection>
<intersection>-217.5 8</intersection>
<intersection>-202 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>434.5,-222.5,437,-222.5</points>
<connection>
<GID>642</GID>
<name>IN_0</name></connection>
<intersection>434.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>434.5,-217.5,437,-217.5</points>
<connection>
<GID>641</GID>
<name>IN_0</name></connection>
<intersection>434.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>287,-135.5,290,-135.5</points>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<connection>
<GID>149</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458.5,-201.5,458.5,-196</points>
<connection>
<GID>640</GID>
<name>SEL_0</name></connection>
<intersection>-196 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432,-196,458.5,-196</points>
<connection>
<GID>644</GID>
<name>IN_0</name></connection>
<intersection>458.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,-138.5,289,-136.5</points>
<intersection>-138.5 1</intersection>
<intersection>-136.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289,-138.5,290,-138.5</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>289 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>287,-136.5,289,-136.5</points>
<connection>
<GID>149</GID>
<name>OUT_2</name></connection>
<intersection>289 0</intersection></hsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455.5,-203,455.5,-199</points>
<intersection>-203 1</intersection>
<intersection>-199 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>455.5,-203,456.5,-203</points>
<connection>
<GID>640</GID>
<name>IN_1</name></connection>
<intersection>455.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>432,-199,455.5,-199</points>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<intersection>455.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,-141.5,288.5,-137.5</points>
<intersection>-141.5 1</intersection>
<intersection>-137.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288.5,-141.5,290,-141.5</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>288.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>287,-137.5,288.5,-137.5</points>
<connection>
<GID>149</GID>
<name>OUT_3</name></connection>
<intersection>288.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>359,-202,376.5,-202</points>
<connection>
<GID>685</GID>
<name>IN_0</name></connection>
<intersection>361.5 5</intersection>
<intersection>376.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>376.5,-204,376.5,-202</points>
<connection>
<GID>661</GID>
<name>IN_0</name></connection>
<intersection>-202 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>361.5,-222.5,361.5,-202</points>
<intersection>-222.5 6</intersection>
<intersection>-217.5 8</intersection>
<intersection>-202 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>361.5,-222.5,364,-222.5</points>
<connection>
<GID>674</GID>
<name>IN_0</name></connection>
<intersection>361.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>361.5,-217.5,364,-217.5</points>
<connection>
<GID>673</GID>
<name>IN_0</name></connection>
<intersection>361.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,-134.5,289,-132.5</points>
<intersection>-134.5 1</intersection>
<intersection>-132.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287,-134.5,289,-134.5</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<intersection>289 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>289,-132.5,290,-132.5</points>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<intersection>289 0</intersection></hsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>460.5,-204,461.5,-204</points>
<connection>
<GID>640</GID>
<name>OUT</name></connection>
<connection>
<GID>653</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>274,-134,279,-134</points>
<connection>
<GID>149</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>152</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>385.5,-201.5,385.5,-196</points>
<connection>
<GID>667</GID>
<name>SEL_0</name></connection>
<intersection>-196 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,-196,385.5,-196</points>
<connection>
<GID>683</GID>
<name>IN_0</name></connection>
<intersection>385.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>382.5,-203,382.5,-199</points>
<intersection>-203 1</intersection>
<intersection>-199 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>382.5,-203,383.5,-203</points>
<connection>
<GID>667</GID>
<name>IN_1</name></connection>
<intersection>382.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>359,-199,382.5,-199</points>
<connection>
<GID>684</GID>
<name>IN_0</name></connection>
<intersection>382.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>387.5,-204,388.5,-204</points>
<connection>
<GID>667</GID>
<name>OUT</name></connection>
<connection>
<GID>688</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382.5,-213,383.5,-213</points>
<connection>
<GID>663</GID>
<name>OUT</name></connection>
<connection>
<GID>689</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>455.5,-213,456.5,-213</points>
<connection>
<GID>635</GID>
<name>OUT</name></connection>
<connection>
<GID>654</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>375,-235.5,377,-235.5</points>
<connection>
<GID>691</GID>
<name>OUT</name></connection>
<connection>
<GID>690</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>377,-251,377,-244.5</points>
<connection>
<GID>692</GID>
<name>IN_2</name></connection>
<intersection>-251 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>375,-251,377,-251</points>
<connection>
<GID>695</GID>
<name>OUT</name></connection>
<intersection>377 0</intersection></hsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>376,-246,376,-242.5</points>
<intersection>-246 2</intersection>
<intersection>-242.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>376,-242.5,377,-242.5</points>
<connection>
<GID>692</GID>
<name>IN_1</name></connection>
<intersection>376 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375,-246,376,-246</points>
<connection>
<GID>694</GID>
<name>OUT</name></connection>
<intersection>376 0</intersection></hsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>375,-240.5,377,-240.5</points>
<connection>
<GID>692</GID>
<name>IN_0</name></connection>
<connection>
<GID>693</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>383,-234.5,384,-234.5</points>
<connection>
<GID>690</GID>
<name>OUT</name></connection>
<connection>
<GID>696</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>360,-234.5,369,-234.5</points>
<connection>
<GID>691</GID>
<name>IN_0</name></connection>
<connection>
<GID>702</GID>
<name>IN_0</name></connection>
<intersection>360 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>360,-245,360,-234.5</points>
<intersection>-245 31</intersection>
<intersection>-239.5 29</intersection>
<intersection>-234.5 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>360,-239.5,369,-239.5</points>
<connection>
<GID>693</GID>
<name>IN_0</name></connection>
<intersection>360 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>360,-245,369,-245</points>
<connection>
<GID>694</GID>
<name>IN_0</name></connection>
<intersection>360 28</intersection></hsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>364,-250,364,-236.5</points>
<intersection>-250 1</intersection>
<intersection>-241.5 4</intersection>
<intersection>-237.5 6</intersection>
<intersection>-236.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>364,-250,369,-250</points>
<connection>
<GID>695</GID>
<name>IN_0</name></connection>
<intersection>364 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>364,-236.5,369,-236.5</points>
<connection>
<GID>691</GID>
<name>IN_1</name></connection>
<intersection>364 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>364,-241.5,369,-241.5</points>
<connection>
<GID>693</GID>
<name>IN_1</name></connection>
<intersection>364 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>360,-237.5,364,-237.5</points>
<connection>
<GID>703</GID>
<name>IN_0</name></connection>
<intersection>364 0</intersection></hsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>368.5,-247,369,-247</points>
<connection>
<GID>697</GID>
<name>OUT_0</name></connection>
<connection>
<GID>694</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>368.5,-252,369,-252</points>
<connection>
<GID>698</GID>
<name>OUT_0</name></connection>
<connection>
<GID>695</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>359.5,-231.5,377,-231.5</points>
<connection>
<GID>701</GID>
<name>IN_0</name></connection>
<intersection>362 5</intersection>
<intersection>377 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>377,-233.5,377,-231.5</points>
<connection>
<GID>690</GID>
<name>IN_0</name></connection>
<intersection>-231.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>362,-252,362,-231.5</points>
<intersection>-252 6</intersection>
<intersection>-247 8</intersection>
<intersection>-231.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>362,-252,364.5,-252</points>
<connection>
<GID>698</GID>
<name>IN_0</name></connection>
<intersection>362 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>362,-247,364.5,-247</points>
<connection>
<GID>697</GID>
<name>IN_0</name></connection>
<intersection>362 5</intersection></hsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>386,-231,386,-225.5</points>
<connection>
<GID>696</GID>
<name>SEL_0</name></connection>
<intersection>-225.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359.5,-225.5,386,-225.5</points>
<connection>
<GID>699</GID>
<name>IN_0</name></connection>
<intersection>386 0</intersection></hsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>383,-232.5,383,-228.5</points>
<intersection>-232.5 1</intersection>
<intersection>-228.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>383,-232.5,384,-232.5</points>
<connection>
<GID>696</GID>
<name>IN_1</name></connection>
<intersection>383 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>359.5,-228.5,383,-228.5</points>
<connection>
<GID>700</GID>
<name>IN_0</name></connection>
<intersection>383 0</intersection></hsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>388,-233.5,389.5,-233.5</points>
<connection>
<GID>696</GID>
<name>OUT</name></connection>
<connection>
<GID>704</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>383,-242.5,384,-242.5</points>
<connection>
<GID>692</GID>
<name>OUT</name></connection>
<connection>
<GID>705</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>448,-235.5,450,-235.5</points>
<connection>
<GID>657</GID>
<name>OUT</name></connection>
<connection>
<GID>656</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>450,-251,450,-244.5</points>
<connection>
<GID>659</GID>
<name>IN_2</name></connection>
<intersection>-251 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>448,-251,450,-251</points>
<connection>
<GID>670</GID>
<name>OUT</name></connection>
<intersection>450 0</intersection></hsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449,-246,449,-242.5</points>
<intersection>-246 2</intersection>
<intersection>-242.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>449,-242.5,450,-242.5</points>
<connection>
<GID>659</GID>
<name>IN_1</name></connection>
<intersection>449 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448,-246,449,-246</points>
<connection>
<GID>669</GID>
<name>OUT</name></connection>
<intersection>449 0</intersection></hsegment></shape></wire>
<wire>
<ID>569</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>448,-240.5,450,-240.5</points>
<connection>
<GID>659</GID>
<name>IN_0</name></connection>
<connection>
<GID>668</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>456,-234.5,457,-234.5</points>
<connection>
<GID>656</GID>
<name>OUT</name></connection>
<connection>
<GID>671</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>433,-234.5,442,-234.5</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<connection>
<GID>679</GID>
<name>IN_0</name></connection>
<intersection>433 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>433,-245,433,-234.5</points>
<intersection>-245 31</intersection>
<intersection>-239.5 29</intersection>
<intersection>-234.5 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>433,-239.5,442,-239.5</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<intersection>433 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>433,-245,442,-245</points>
<connection>
<GID>669</GID>
<name>IN_0</name></connection>
<intersection>433 28</intersection></hsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>437,-250,437,-236.5</points>
<intersection>-250 1</intersection>
<intersection>-241.5 4</intersection>
<intersection>-237.5 6</intersection>
<intersection>-236.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>437,-250,442,-250</points>
<connection>
<GID>670</GID>
<name>IN_0</name></connection>
<intersection>437 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>437,-236.5,442,-236.5</points>
<connection>
<GID>657</GID>
<name>IN_1</name></connection>
<intersection>437 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>437,-241.5,442,-241.5</points>
<connection>
<GID>668</GID>
<name>IN_1</name></connection>
<intersection>437 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>433,-237.5,437,-237.5</points>
<connection>
<GID>680</GID>
<name>IN_0</name></connection>
<intersection>437 0</intersection></hsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>441.5,-247,442,-247</points>
<connection>
<GID>672</GID>
<name>OUT_0</name></connection>
<connection>
<GID>669</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>574</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>441.5,-252,442,-252</points>
<connection>
<GID>675</GID>
<name>OUT_0</name></connection>
<connection>
<GID>670</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432.5,-231.5,450,-231.5</points>
<connection>
<GID>678</GID>
<name>IN_0</name></connection>
<intersection>435 5</intersection>
<intersection>450 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>450,-233.5,450,-231.5</points>
<connection>
<GID>656</GID>
<name>IN_0</name></connection>
<intersection>-231.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>435,-252,435,-231.5</points>
<intersection>-252 6</intersection>
<intersection>-247 8</intersection>
<intersection>-231.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>435,-252,437.5,-252</points>
<connection>
<GID>675</GID>
<name>IN_0</name></connection>
<intersection>435 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>435,-247,437.5,-247</points>
<connection>
<GID>672</GID>
<name>IN_0</name></connection>
<intersection>435 5</intersection></hsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459,-231,459,-225.5</points>
<connection>
<GID>671</GID>
<name>SEL_0</name></connection>
<intersection>-225.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432.5,-225.5,459,-225.5</points>
<connection>
<GID>676</GID>
<name>IN_0</name></connection>
<intersection>459 0</intersection></hsegment></shape></wire>
<wire>
<ID>577</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,-232.5,456,-228.5</points>
<intersection>-232.5 1</intersection>
<intersection>-228.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>456,-232.5,457,-232.5</points>
<connection>
<GID>671</GID>
<name>IN_1</name></connection>
<intersection>456 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>432.5,-228.5,456,-228.5</points>
<connection>
<GID>677</GID>
<name>IN_0</name></connection>
<intersection>456 0</intersection></hsegment></shape></wire>
<wire>
<ID>578</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>461,-233.5,462.5,-233.5</points>
<connection>
<GID>671</GID>
<name>OUT</name></connection>
<connection>
<GID>681</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>579</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>456,-242.5,457,-242.5</points>
<connection>
<GID>659</GID>
<name>OUT</name></connection>
<connection>
<GID>682</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>580</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>457,-304,467,-304</points>
<connection>
<GID>596</GID>
<name>OUT</name></connection>
<connection>
<GID>707</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>581</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-158,278,-151.5</points>
<intersection>-158 2</intersection>
<intersection>-151.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274,-151.5,278,-151.5</points>
<connection>
<GID>709</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>278,-158,279,-158</points>
<connection>
<GID>613</GID>
<name>IN_B_0</name></connection>
<intersection>278 0</intersection></hsegment></shape></wire>
<wire>
<ID>582</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>274,-165,279,-165</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<connection>
<GID>623</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-168.5,276,-166</points>
<intersection>-168.5 2</intersection>
<intersection>-166 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-166,279,-166</points>
<connection>
<GID>613</GID>
<name>IN_1</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274,-168.5,276,-168.5</points>
<connection>
<GID>625</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>584</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277,-171.5,277,-167</points>
<intersection>-171.5 2</intersection>
<intersection>-167 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277,-167,279,-167</points>
<connection>
<GID>613</GID>
<name>IN_2</name></connection>
<intersection>277 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274,-171.5,277,-171.5</points>
<connection>
<GID>627</GID>
<name>IN_0</name></connection>
<intersection>277 0</intersection></hsegment></shape></wire>
<wire>
<ID>585</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-174.5,278,-168</points>
<intersection>-174.5 2</intersection>
<intersection>-168 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>278,-168,279,-168</points>
<connection>
<GID>613</GID>
<name>IN_3</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274,-174.5,278,-174.5</points>
<connection>
<GID>631</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment></shape></wire>
<wire>
<ID>586</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>287,-189.5,290,-189.5</points>
<connection>
<GID>711</GID>
<name>IN_0</name></connection>
<connection>
<GID>714</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>587</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,-192.5,289,-190.5</points>
<intersection>-192.5 1</intersection>
<intersection>-190.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289,-192.5,290,-192.5</points>
<connection>
<GID>712</GID>
<name>IN_0</name></connection>
<intersection>289 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>287,-190.5,289,-190.5</points>
<connection>
<GID>714</GID>
<name>OUT_2</name></connection>
<intersection>289 0</intersection></hsegment></shape></wire>
<wire>
<ID>588</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,-195.5,288.5,-191.5</points>
<intersection>-195.5 1</intersection>
<intersection>-191.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288.5,-195.5,290,-195.5</points>
<connection>
<GID>713</GID>
<name>IN_0</name></connection>
<intersection>288.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>287,-191.5,288.5,-191.5</points>
<connection>
<GID>714</GID>
<name>OUT_3</name></connection>
<intersection>288.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,-188.5,289,-186.5</points>
<intersection>-188.5 1</intersection>
<intersection>-186.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287,-188.5,289,-188.5</points>
<connection>
<GID>714</GID>
<name>OUT_0</name></connection>
<intersection>289 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>289,-186.5,290,-186.5</points>
<connection>
<GID>710</GID>
<name>IN_0</name></connection>
<intersection>289 0</intersection></hsegment></shape></wire>
<wire>
<ID>590</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>274,-188,279,-188</points>
<connection>
<GID>714</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>715</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-133,276,-130.5</points>
<intersection>-133 2</intersection>
<intersection>-130.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274,-130.5,276,-130.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-133,279,-133</points>
<connection>
<GID>149</GID>
<name>IN_B_2</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-187,276,-184.5</points>
<intersection>-187 2</intersection>
<intersection>-184.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274,-184.5,276,-184.5</points>
<connection>
<GID>720</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-187,279,-187</points>
<connection>
<GID>714</GID>
<name>IN_B_2</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277,-132,277,-127.5</points>
<intersection>-132 2</intersection>
<intersection>-127.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274,-127.5,277,-127.5</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>277 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277,-132,279,-132</points>
<connection>
<GID>149</GID>
<name>IN_B_1</name></connection>
<intersection>277 0</intersection></hsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277,-186,277,-181.5</points>
<intersection>-186 2</intersection>
<intersection>-181.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274.5,-181.5,277,-181.5</points>
<connection>
<GID>721</GID>
<name>IN_0</name></connection>
<intersection>277 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277,-186,279,-186</points>
<connection>
<GID>714</GID>
<name>IN_B_1</name></connection>
<intersection>277 0</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-131,278,-124.5</points>
<intersection>-131 2</intersection>
<intersection>-124.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274,-124.5,278,-124.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>278,-131,279,-131</points>
<connection>
<GID>149</GID>
<name>IN_B_0</name></connection>
<intersection>278 0</intersection></hsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-185,278,-178.5</points>
<intersection>-185 2</intersection>
<intersection>-178.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274,-178.5,278,-178.5</points>
<connection>
<GID>722</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>278,-185,279,-185</points>
<connection>
<GID>714</GID>
<name>IN_B_0</name></connection>
<intersection>278 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>374,-141,376,-141</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<connection>
<GID>301</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>274,-192,279,-192</points>
<connection>
<GID>714</GID>
<name>IN_0</name></connection>
<connection>
<GID>716</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>376,-156.5,376,-150</points>
<connection>
<GID>303</GID>
<name>IN_2</name></connection>
<intersection>-156.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>374,-156.5,376,-156.5</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<intersection>376 0</intersection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-195.5,276,-193</points>
<intersection>-195.5 2</intersection>
<intersection>-193 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-193,279,-193</points>
<connection>
<GID>714</GID>
<name>IN_1</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274,-195.5,276,-195.5</points>
<connection>
<GID>717</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375,-151.5,375,-148</points>
<intersection>-151.5 2</intersection>
<intersection>-148 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375,-148,376,-148</points>
<connection>
<GID>303</GID>
<name>IN_1</name></connection>
<intersection>375 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>374,-151.5,375,-151.5</points>
<connection>
<GID>313</GID>
<name>OUT</name></connection>
<intersection>375 0</intersection></hsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277,-198.5,277,-194</points>
<intersection>-198.5 2</intersection>
<intersection>-194 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277,-194,279,-194</points>
<connection>
<GID>714</GID>
<name>IN_2</name></connection>
<intersection>277 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274,-198.5,277,-198.5</points>
<connection>
<GID>718</GID>
<name>IN_0</name></connection>
<intersection>277 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>374,-146,376,-146</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<connection>
<GID>309</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-201.5,278,-195</points>
<intersection>-201.5 2</intersection>
<intersection>-195 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>278,-195,279,-195</points>
<connection>
<GID>714</GID>
<name>IN_3</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274,-201.5,278,-201.5</points>
<connection>
<GID>719</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>287,-216.5,290,-216.5</points>
<connection>
<GID>724</GID>
<name>IN_0</name></connection>
<connection>
<GID>727</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,-219.5,289,-217.5</points>
<intersection>-219.5 1</intersection>
<intersection>-217.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289,-219.5,290,-219.5</points>
<connection>
<GID>725</GID>
<name>IN_0</name></connection>
<intersection>289 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>287,-217.5,289,-217.5</points>
<connection>
<GID>727</GID>
<name>OUT_2</name></connection>
<intersection>289 0</intersection></hsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,-222.5,288.5,-218.5</points>
<intersection>-222.5 1</intersection>
<intersection>-218.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288.5,-222.5,290,-222.5</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<intersection>288.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>287,-218.5,288.5,-218.5</points>
<connection>
<GID>727</GID>
<name>OUT_3</name></connection>
<intersection>288.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382,-140,383,-140</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<connection>
<GID>301</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,-215.5,289,-213.5</points>
<intersection>-215.5 1</intersection>
<intersection>-213.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287,-215.5,289,-215.5</points>
<connection>
<GID>727</GID>
<name>OUT_0</name></connection>
<intersection>289 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>289,-213.5,290,-213.5</points>
<connection>
<GID>723</GID>
<name>IN_0</name></connection>
<intersection>289 0</intersection></hsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>274,-215,279,-215</points>
<connection>
<GID>727</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>728</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>359,-140,368,-140</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<intersection>365.5 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>365.5,-150.5,365.5,-140</points>
<intersection>-150.5 31</intersection>
<intersection>-145 29</intersection>
<intersection>-140 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>365.5,-145,368,-145</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>365.5 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>365.5,-150.5,368,-150.5</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>365.5 28</intersection></hsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-214,276,-211.5</points>
<intersection>-214 2</intersection>
<intersection>-211.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274,-211.5,276,-211.5</points>
<connection>
<GID>733</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-214,279,-214</points>
<connection>
<GID>727</GID>
<name>IN_B_2</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363,-155.5,363,-142</points>
<intersection>-155.5 1</intersection>
<intersection>-147 4</intersection>
<intersection>-143 6</intersection>
<intersection>-142 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>363,-155.5,368,-155.5</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>363 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>363,-142,368,-142</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>363 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>363,-147,368,-147</points>
<connection>
<GID>309</GID>
<name>IN_1</name></connection>
<intersection>363 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>359,-143,363,-143</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>363 0</intersection></hsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277,-213,277,-208.5</points>
<intersection>-213 2</intersection>
<intersection>-208.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274,-208.5,277,-208.5</points>
<connection>
<GID>734</GID>
<name>IN_0</name></connection>
<intersection>277 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277,-213,279,-213</points>
<connection>
<GID>727</GID>
<name>IN_B_1</name></connection>
<intersection>277 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>367.5,-152.5,368,-152.5</points>
<connection>
<GID>316</GID>
<name>OUT_0</name></connection>
<connection>
<GID>313</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-212,278,-205.5</points>
<intersection>-212 2</intersection>
<intersection>-205.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274,-205.5,278,-205.5</points>
<connection>
<GID>735</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>278,-212,279,-212</points>
<connection>
<GID>727</GID>
<name>IN_B_0</name></connection>
<intersection>278 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>367.5,-157.5,368,-157.5</points>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection>
<connection>
<GID>314</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>274,-219,279,-219</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<connection>
<GID>729</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-222.5,276,-220</points>
<intersection>-222.5 2</intersection>
<intersection>-220 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-220,279,-220</points>
<connection>
<GID>727</GID>
<name>IN_1</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274,-222.5,276,-222.5</points>
<connection>
<GID>730</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>358.5,-137,376,-137</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>361 5</intersection>
<intersection>376 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>376,-139,376,-137</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>-137 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>361,-157.5,361,-137</points>
<intersection>-157.5 6</intersection>
<intersection>-152.5 8</intersection>
<intersection>-137 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>361,-157.5,363.5,-157.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>361 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>361,-152.5,363.5,-152.5</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>361 5</intersection></hsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277,-225.5,277,-221</points>
<intersection>-225.5 2</intersection>
<intersection>-221 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277,-221,279,-221</points>
<connection>
<GID>727</GID>
<name>IN_2</name></connection>
<intersection>277 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274,-225.5,277,-225.5</points>
<connection>
<GID>731</GID>
<name>IN_0</name></connection>
<intersection>277 0</intersection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-228.5,278,-222</points>
<intersection>-228.5 2</intersection>
<intersection>-222 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>278,-222,279,-222</points>
<connection>
<GID>727</GID>
<name>IN_3</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274,-228.5,278,-228.5</points>
<connection>
<GID>732</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-155,282,-144</points>
<connection>
<GID>149</GID>
<name>carry_out</name></connection>
<connection>
<GID>613</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-182,282,-171</points>
<connection>
<GID>613</GID>
<name>carry_out</name></connection>
<connection>
<GID>714</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-209,282,-198</points>
<connection>
<GID>714</GID>
<name>carry_out</name></connection>
<connection>
<GID>727</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>385,-136.5,385,-131</points>
<connection>
<GID>315</GID>
<name>SEL_0</name></connection>
<intersection>-131 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>358.5,-131,385,-131</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>385 0</intersection></hsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-128,282,-124.5</points>
<connection>
<GID>149</GID>
<name>carry_in</name></connection>
<intersection>-124.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>285,-126,285,-124.5</points>
<connection>
<GID>737</GID>
<name>OUT_0</name></connection>
<intersection>-124.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>282,-124.5,285,-124.5</points>
<intersection>282 0</intersection>
<intersection>285 1</intersection></hsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-228,282,-225</points>
<connection>
<GID>727</GID>
<name>carry_out</name></connection>
<intersection>-228 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282,-228,299.5,-228</points>
<connection>
<GID>739</GID>
<name>N_in0</name></connection>
<intersection>282 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>382,-138,382,-134</points>
<intersection>-138 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>382,-138,383,-138</points>
<connection>
<GID>315</GID>
<name>IN_1</name></connection>
<intersection>382 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>358.5,-134,382,-134</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>382 0</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>387,-139,388,-139</points>
<connection>
<GID>315</GID>
<name>OUT</name></connection>
<connection>
<GID>418</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382,-148,383,-148</points>
<connection>
<GID>303</GID>
<name>OUT</name></connection>
<connection>
<GID>419</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>374.5,-170.5,376.5,-170.5</points>
<connection>
<GID>423</GID>
<name>OUT</name></connection>
<connection>
<GID>421</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>376.5,-186,376.5,-179.5</points>
<connection>
<GID>425</GID>
<name>IN_2</name></connection>
<intersection>-186 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>374.5,-186,376.5,-186</points>
<connection>
<GID>435</GID>
<name>OUT</name></connection>
<intersection>376.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375.5,-181,375.5,-177.5</points>
<intersection>-181 2</intersection>
<intersection>-177.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375.5,-177.5,376.5,-177.5</points>
<connection>
<GID>425</GID>
<name>IN_1</name></connection>
<intersection>375.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>374.5,-181,375.5,-181</points>
<connection>
<GID>429</GID>
<name>OUT</name></connection>
<intersection>375.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>374,-175.5,376.5,-175.5</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<connection>
<GID>427</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382.5,-169.5,383.5,-169.5</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<connection>
<GID>421</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>359.5,-169.5,368.5,-169.5</points>
<connection>
<GID>423</GID>
<name>IN_0</name></connection>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>366 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>366,-180,366,-169.5</points>
<intersection>-180 31</intersection>
<intersection>-174.5 29</intersection>
<intersection>-169.5 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>366,-174.5,368,-174.5</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<intersection>366 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>366,-180,368.5,-180</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<intersection>366 28</intersection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363.5,-185,363.5,-171.5</points>
<intersection>-185 1</intersection>
<intersection>-176.5 4</intersection>
<intersection>-172.5 6</intersection>
<intersection>-171.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>363.5,-185,368.5,-185</points>
<connection>
<GID>435</GID>
<name>IN_0</name></connection>
<intersection>363.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>363.5,-171.5,368.5,-171.5</points>
<connection>
<GID>423</GID>
<name>IN_1</name></connection>
<intersection>363.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>363.5,-176.5,368,-176.5</points>
<connection>
<GID>427</GID>
<name>IN_1</name></connection>
<intersection>363.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>359.5,-172.5,363.5,-172.5</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>363.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>368,-182,368.5,-182</points>
<connection>
<GID>437</GID>
<name>OUT_0</name></connection>
<connection>
<GID>429</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>368,-187,368.5,-187</points>
<connection>
<GID>438</GID>
<name>OUT_0</name></connection>
<connection>
<GID>435</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>359,-166.5,376.5,-166.5</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<intersection>361.5 5</intersection>
<intersection>376.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>376.5,-168.5,376.5,-166.5</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<intersection>-166.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>361.5,-187,361.5,-166.5</points>
<intersection>-187 6</intersection>
<intersection>-182 8</intersection>
<intersection>-166.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>361.5,-187,364,-187</points>
<connection>
<GID>438</GID>
<name>IN_0</name></connection>
<intersection>361.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>361.5,-182,364,-182</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<intersection>361.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>385.5,-166,385.5,-160.5</points>
<connection>
<GID>436</GID>
<name>SEL_0</name></connection>
<intersection>-160.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,-160.5,385.5,-160.5</points>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<intersection>385.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>382.5,-167.5,382.5,-163.5</points>
<intersection>-167.5 1</intersection>
<intersection>-163.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>382.5,-167.5,383.5,-167.5</points>
<connection>
<GID>436</GID>
<name>IN_1</name></connection>
<intersection>382.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>359,-163.5,382.5,-163.5</points>
<connection>
<GID>440</GID>
<name>IN_0</name></connection>
<intersection>382.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>387.5,-168.5,389.5,-168.5</points>
<connection>
<GID>436</GID>
<name>OUT</name></connection>
<connection>
<GID>453</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382.5,-177.5,383.5,-177.5</points>
<connection>
<GID>425</GID>
<name>OUT</name></connection>
<connection>
<GID>455</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>274,-138,279,-138</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<connection>
<GID>158</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>447,-141,449,-141</points>
<connection>
<GID>484</GID>
<name>OUT</name></connection>
<connection>
<GID>482</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449,-156.5,449,-150</points>
<connection>
<GID>485</GID>
<name>IN_2</name></connection>
<intersection>-156.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>447,-156.5,449,-156.5</points>
<connection>
<GID>489</GID>
<name>OUT</name></connection>
<intersection>449 0</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448,-151.5,448,-148</points>
<intersection>-151.5 2</intersection>
<intersection>-148 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>448,-148,449,-148</points>
<connection>
<GID>485</GID>
<name>IN_1</name></connection>
<intersection>448 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447,-151.5,448,-151.5</points>
<connection>
<GID>488</GID>
<name>OUT</name></connection>
<intersection>448 0</intersection></hsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>447,-146,449,-146</points>
<connection>
<GID>485</GID>
<name>IN_0</name></connection>
<connection>
<GID>487</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>455,-140,456,-140</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<connection>
<GID>482</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432,-140,441,-140</points>
<connection>
<GID>484</GID>
<name>IN_0</name></connection>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<intersection>438.5 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>438.5,-150.5,438.5,-140</points>
<intersection>-150.5 31</intersection>
<intersection>-145 29</intersection>
<intersection>-140 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>438.5,-145,441,-145</points>
<connection>
<GID>487</GID>
<name>IN_0</name></connection>
<intersection>438.5 28</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>438.5,-150.5,441,-150.5</points>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<intersection>438.5 28</intersection></hsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-141.5,276,-139</points>
<intersection>-141.5 2</intersection>
<intersection>-139 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-139,279,-139</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274,-141.5,276,-141.5</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277,-144.5,277,-140</points>
<intersection>-144.5 2</intersection>
<intersection>-140 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277,-140,279,-140</points>
<connection>
<GID>149</GID>
<name>IN_2</name></connection>
<intersection>277 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274,-144.5,277,-144.5</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>277 0</intersection></hsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-147,278,-141</points>
<intersection>-147 2</intersection>
<intersection>-141 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>278,-141,279,-141</points>
<connection>
<GID>149</GID>
<name>IN_3</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274,-147,278,-147</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>287,-162.5,290,-162.5</points>
<connection>
<GID>609</GID>
<name>IN_0</name></connection>
<connection>
<GID>613</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436,-155.5,436,-142</points>
<intersection>-155.5 1</intersection>
<intersection>-147 4</intersection>
<intersection>-143 6</intersection>
<intersection>-142 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>436,-155.5,441,-155.5</points>
<connection>
<GID>489</GID>
<name>IN_0</name></connection>
<intersection>436 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>436,-142,441,-142</points>
<connection>
<GID>484</GID>
<name>IN_1</name></connection>
<intersection>436 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>436,-147,441,-147</points>
<connection>
<GID>487</GID>
<name>IN_1</name></connection>
<intersection>436 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>432,-143,436,-143</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>436 0</intersection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440.5,-152.5,441,-152.5</points>
<connection>
<GID>491</GID>
<name>OUT_0</name></connection>
<connection>
<GID>488</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>386</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440.5,-157.5,441,-157.5</points>
<connection>
<GID>492</GID>
<name>OUT_0</name></connection>
<connection>
<GID>489</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>431.5,-137,449,-137</points>
<connection>
<GID>497</GID>
<name>IN_0</name></connection>
<intersection>434 5</intersection>
<intersection>449 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>449,-139,449,-137</points>
<connection>
<GID>482</GID>
<name>IN_0</name></connection>
<intersection>-137 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>434,-157.5,434,-137</points>
<intersection>-157.5 6</intersection>
<intersection>-152.5 8</intersection>
<intersection>-137 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>434,-157.5,436.5,-157.5</points>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<intersection>434 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>434,-152.5,436.5,-152.5</points>
<connection>
<GID>491</GID>
<name>IN_0</name></connection>
<intersection>434 5</intersection></hsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458,-136.5,458,-131</points>
<connection>
<GID>490</GID>
<name>SEL_0</name></connection>
<intersection>-131 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>431.5,-131,458,-131</points>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<intersection>458 0</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>636.148,49.6298,1133.01,-206.626</PageViewport>
<gate>
<ID>772</ID>
<type>DA_FROM</type>
<position>652,-42</position>
<input>
<ID>IN_0</ID>636 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_RAM</lparam></gate>
<gate>
<ID>773</ID>
<type>DE_TO</type>
<position>662,-40</position>
<input>
<ID>IN_0</ID>637 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_MUX_OUT</lparam></gate>
<gate>
<ID>774</ID>
<type>DA_FROM</type>
<position>652,-36</position>
<input>
<ID>IN_0</ID>638 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>775</ID>
<type>AA_MUX_2x1</type>
<position>657,-49</position>
<input>
<ID>IN_0</ID>640 </input>
<input>
<ID>IN_1</ID>639 </input>
<output>
<ID>OUT</ID>641 </output>
<input>
<ID>SEL_0</ID>642 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>776</ID>
<type>DA_FROM</type>
<position>652,-48</position>
<input>
<ID>IN_0</ID>639 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_ES</lparam></gate>
<gate>
<ID>777</ID>
<type>DA_FROM</type>
<position>652,-51</position>
<input>
<ID>IN_0</ID>640 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_RAM</lparam></gate>
<gate>
<ID>778</ID>
<type>DE_TO</type>
<position>662,-49</position>
<input>
<ID>IN_0</ID>641 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6_MUX_OUT</lparam></gate>
<gate>
<ID>779</ID>
<type>DA_FROM</type>
<position>652,-45</position>
<input>
<ID>IN_0</ID>642 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>780</ID>
<type>AA_MUX_2x1</type>
<position>657,-58</position>
<input>
<ID>IN_0</ID>644 </input>
<input>
<ID>IN_1</ID>643 </input>
<output>
<ID>OUT</ID>645 </output>
<input>
<ID>SEL_0</ID>646 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>781</ID>
<type>DA_FROM</type>
<position>652,-57</position>
<input>
<ID>IN_0</ID>643 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_ES</lparam></gate>
<gate>
<ID>782</ID>
<type>DA_FROM</type>
<position>652,-60</position>
<input>
<ID>IN_0</ID>644 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_RAM</lparam></gate>
<gate>
<ID>783</ID>
<type>DE_TO</type>
<position>662,-58</position>
<input>
<ID>IN_0</ID>645 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7_MUX_OUT</lparam></gate>
<gate>
<ID>784</ID>
<type>DA_FROM</type>
<position>652,-54</position>
<input>
<ID>IN_0</ID>646 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>785</ID>
<type>AA_MUX_2x1</type>
<position>717,5.5</position>
<input>
<ID>IN_0</ID>648 </input>
<input>
<ID>IN_1</ID>647 </input>
<output>
<ID>OUT</ID>649 </output>
<input>
<ID>SEL_0</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>786</ID>
<type>DA_FROM</type>
<position>712,6.5</position>
<input>
<ID>IN_0</ID>647 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_ES</lparam></gate>
<gate>
<ID>787</ID>
<type>DA_FROM</type>
<position>712,3.5</position>
<input>
<ID>IN_0</ID>648 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_RAM</lparam></gate>
<gate>
<ID>788</ID>
<type>DE_TO</type>
<position>722,5.5</position>
<input>
<ID>IN_0</ID>649 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8_MUX_OUT</lparam></gate>
<gate>
<ID>789</ID>
<type>DA_FROM</type>
<position>712,9.5</position>
<input>
<ID>IN_0</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>790</ID>
<type>AA_MUX_2x1</type>
<position>717,-3.5</position>
<input>
<ID>IN_0</ID>652 </input>
<input>
<ID>IN_1</ID>651 </input>
<output>
<ID>OUT</ID>653 </output>
<input>
<ID>SEL_0</ID>654 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>791</ID>
<type>DA_FROM</type>
<position>712,-2.5</position>
<input>
<ID>IN_0</ID>651 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_ES</lparam></gate>
<gate>
<ID>792</ID>
<type>DA_FROM</type>
<position>712,-5.5</position>
<input>
<ID>IN_0</ID>652 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_RAM</lparam></gate>
<gate>
<ID>793</ID>
<type>DE_TO</type>
<position>722,-3.5</position>
<input>
<ID>IN_0</ID>653 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9_MUX_OUT</lparam></gate>
<gate>
<ID>794</ID>
<type>DA_FROM</type>
<position>712,0.5</position>
<input>
<ID>IN_0</ID>654 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>795</ID>
<type>AA_MUX_2x1</type>
<position>717,-12.5</position>
<input>
<ID>IN_0</ID>656 </input>
<input>
<ID>IN_1</ID>655 </input>
<output>
<ID>OUT</ID>657 </output>
<input>
<ID>SEL_0</ID>658 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>796</ID>
<type>DA_FROM</type>
<position>712,-11.5</position>
<input>
<ID>IN_0</ID>655 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_ES</lparam></gate>
<gate>
<ID>797</ID>
<type>DA_FROM</type>
<position>712,-14.5</position>
<input>
<ID>IN_0</ID>656 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_RAM</lparam></gate>
<gate>
<ID>798</ID>
<type>DE_TO</type>
<position>722,-12.5</position>
<input>
<ID>IN_0</ID>657 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10_MUX_OUT</lparam></gate>
<gate>
<ID>799</ID>
<type>DA_FROM</type>
<position>712,-8.5</position>
<input>
<ID>IN_0</ID>658 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>800</ID>
<type>AA_MUX_2x1</type>
<position>717,-21.5</position>
<input>
<ID>IN_0</ID>660 </input>
<input>
<ID>IN_1</ID>659 </input>
<output>
<ID>OUT</ID>661 </output>
<input>
<ID>SEL_0</ID>662 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>801</ID>
<type>DA_FROM</type>
<position>712,-20.5</position>
<input>
<ID>IN_0</ID>659 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_ES</lparam></gate>
<gate>
<ID>802</ID>
<type>DA_FROM</type>
<position>712,-23.5</position>
<input>
<ID>IN_0</ID>660 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_RAM</lparam></gate>
<gate>
<ID>803</ID>
<type>DE_TO</type>
<position>722,-21.5</position>
<input>
<ID>IN_0</ID>661 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11_MUX_OUT</lparam></gate>
<gate>
<ID>804</ID>
<type>DA_FROM</type>
<position>712,-17.5</position>
<input>
<ID>IN_0</ID>662 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>805</ID>
<type>AA_MUX_2x1</type>
<position>717,-30.5</position>
<input>
<ID>IN_0</ID>664 </input>
<input>
<ID>IN_1</ID>663 </input>
<output>
<ID>OUT</ID>665 </output>
<input>
<ID>SEL_0</ID>666 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>806</ID>
<type>DA_FROM</type>
<position>712,-29.5</position>
<input>
<ID>IN_0</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_ES</lparam></gate>
<gate>
<ID>807</ID>
<type>DA_FROM</type>
<position>712,-32.5</position>
<input>
<ID>IN_0</ID>664 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_RAM</lparam></gate>
<gate>
<ID>808</ID>
<type>DE_TO</type>
<position>722,-30.5</position>
<input>
<ID>IN_0</ID>665 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_MUX_OUT</lparam></gate>
<gate>
<ID>809</ID>
<type>DA_FROM</type>
<position>712,-26.5</position>
<input>
<ID>IN_0</ID>666 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>810</ID>
<type>AA_MUX_2x1</type>
<position>717,-39.5</position>
<input>
<ID>IN_0</ID>668 </input>
<input>
<ID>IN_1</ID>667 </input>
<output>
<ID>OUT</ID>669 </output>
<input>
<ID>SEL_0</ID>670 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>811</ID>
<type>DA_FROM</type>
<position>712,-38.5</position>
<input>
<ID>IN_0</ID>667 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_ES</lparam></gate>
<gate>
<ID>812</ID>
<type>DA_FROM</type>
<position>712,-41.5</position>
<input>
<ID>IN_0</ID>668 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_RAM</lparam></gate>
<gate>
<ID>813</ID>
<type>DE_TO</type>
<position>722,-39.5</position>
<input>
<ID>IN_0</ID>669 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_MUX_OUT</lparam></gate>
<gate>
<ID>814</ID>
<type>DA_FROM</type>
<position>712,-35.5</position>
<input>
<ID>IN_0</ID>670 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>815</ID>
<type>AA_MUX_2x1</type>
<position>717,-48.5</position>
<input>
<ID>IN_0</ID>672 </input>
<input>
<ID>IN_1</ID>671 </input>
<output>
<ID>OUT</ID>673 </output>
<input>
<ID>SEL_0</ID>674 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>816</ID>
<type>DA_FROM</type>
<position>712,-47.5</position>
<input>
<ID>IN_0</ID>671 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_ES</lparam></gate>
<gate>
<ID>817</ID>
<type>DA_FROM</type>
<position>712,-50.5</position>
<input>
<ID>IN_0</ID>672 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_RAM</lparam></gate>
<gate>
<ID>818</ID>
<type>DE_TO</type>
<position>722,-48.5</position>
<input>
<ID>IN_0</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_MUX_OUT</lparam></gate>
<gate>
<ID>819</ID>
<type>DA_FROM</type>
<position>712,-44.5</position>
<input>
<ID>IN_0</ID>674 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>820</ID>
<type>AA_MUX_2x1</type>
<position>717,-57.5</position>
<input>
<ID>IN_0</ID>676 </input>
<input>
<ID>IN_1</ID>675 </input>
<output>
<ID>OUT</ID>677 </output>
<input>
<ID>SEL_0</ID>678 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>821</ID>
<type>DA_FROM</type>
<position>712,-56.5</position>
<input>
<ID>IN_0</ID>675 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_ES</lparam></gate>
<gate>
<ID>822</ID>
<type>DA_FROM</type>
<position>712,-59.5</position>
<input>
<ID>IN_0</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_RAM</lparam></gate>
<gate>
<ID>823</ID>
<type>DE_TO</type>
<position>722,-57.5</position>
<input>
<ID>IN_0</ID>677 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_MUX_OUT</lparam></gate>
<gate>
<ID>824</ID>
<type>DA_FROM</type>
<position>712,-53.5</position>
<input>
<ID>IN_0</ID>678 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>826</ID>
<type>AA_LABEL</type>
<position>685.5,16</position>
<gparam>LABEL_TEXT Mux</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>263</ID>
<type>AA_LABEL</type>
<position>666,26</position>
<gparam>LABEL_TEXT Prof.  Angelo Zanini / Nuncio Perrella</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>266</ID>
<type>AA_LABEL</type>
<position>674.5,34</position>
<gparam>LABEL_TEXT PROCESSADOR BIP IMT - MAUA 2022</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>871</ID>
<type>AA_LABEL</type>
<position>591.5,-6.5</position>
<gparam>LABEL_TEXT Sinais de Controle</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>872</ID>
<type>AA_LABEL</type>
<position>588.5,-15</position>
<gparam>LABEL_TEXT SelUlaSrc</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>741</ID>
<type>AA_MUX_2x1</type>
<position>657,6</position>
<input>
<ID>IN_0</ID>616 </input>
<input>
<ID>IN_1</ID>615 </input>
<output>
<ID>OUT</ID>617 </output>
<input>
<ID>SEL_0</ID>618 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>743</ID>
<type>DA_FROM</type>
<position>652,7</position>
<input>
<ID>IN_0</ID>615 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_ES</lparam></gate>
<gate>
<ID>745</ID>
<type>DA_FROM</type>
<position>652,4</position>
<input>
<ID>IN_0</ID>616 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_RAM</lparam></gate>
<gate>
<ID>747</ID>
<type>DE_TO</type>
<position>662,6</position>
<input>
<ID>IN_0</ID>617 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0_MUX_OUT</lparam></gate>
<gate>
<ID>749</ID>
<type>DA_FROM</type>
<position>652,10</position>
<input>
<ID>IN_0</ID>618 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>750</ID>
<type>AA_MUX_2x1</type>
<position>657,-4</position>
<input>
<ID>IN_0</ID>620 </input>
<input>
<ID>IN_1</ID>619 </input>
<output>
<ID>OUT</ID>621 </output>
<input>
<ID>SEL_0</ID>622 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>751</ID>
<type>DA_FROM</type>
<position>652,-3</position>
<input>
<ID>IN_0</ID>619 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_ES</lparam></gate>
<gate>
<ID>752</ID>
<type>DA_FROM</type>
<position>652,-6</position>
<input>
<ID>IN_0</ID>620 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_RAM</lparam></gate>
<gate>
<ID>753</ID>
<type>DE_TO</type>
<position>662,-4</position>
<input>
<ID>IN_0</ID>621 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1_MUX_OUT</lparam></gate>
<gate>
<ID>754</ID>
<type>DA_FROM</type>
<position>652,0</position>
<input>
<ID>IN_0</ID>622 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>755</ID>
<type>AA_MUX_2x1</type>
<position>657,-13</position>
<input>
<ID>IN_0</ID>624 </input>
<input>
<ID>IN_1</ID>623 </input>
<output>
<ID>OUT</ID>625 </output>
<input>
<ID>SEL_0</ID>626 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>756</ID>
<type>DA_FROM</type>
<position>652,-12</position>
<input>
<ID>IN_0</ID>623 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_ES</lparam></gate>
<gate>
<ID>757</ID>
<type>DA_FROM</type>
<position>652,-15</position>
<input>
<ID>IN_0</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_RAM</lparam></gate>
<gate>
<ID>758</ID>
<type>DE_TO</type>
<position>662,-13</position>
<input>
<ID>IN_0</ID>625 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2_MUX_OUT</lparam></gate>
<gate>
<ID>759</ID>
<type>DA_FROM</type>
<position>652,-9</position>
<input>
<ID>IN_0</ID>626 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>760</ID>
<type>AA_MUX_2x1</type>
<position>657,-22</position>
<input>
<ID>IN_0</ID>628 </input>
<input>
<ID>IN_1</ID>627 </input>
<output>
<ID>OUT</ID>629 </output>
<input>
<ID>SEL_0</ID>630 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>761</ID>
<type>DA_FROM</type>
<position>652,-21</position>
<input>
<ID>IN_0</ID>627 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_ES</lparam></gate>
<gate>
<ID>762</ID>
<type>DA_FROM</type>
<position>652,-24</position>
<input>
<ID>IN_0</ID>628 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_RAM</lparam></gate>
<gate>
<ID>763</ID>
<type>DE_TO</type>
<position>662,-22</position>
<input>
<ID>IN_0</ID>629 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3_MUX_OUT</lparam></gate>
<gate>
<ID>764</ID>
<type>DA_FROM</type>
<position>652,-18</position>
<input>
<ID>IN_0</ID>630 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>765</ID>
<type>AA_MUX_2x1</type>
<position>657,-31</position>
<input>
<ID>IN_0</ID>632 </input>
<input>
<ID>IN_1</ID>631 </input>
<output>
<ID>OUT</ID>633 </output>
<input>
<ID>SEL_0</ID>634 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>766</ID>
<type>DA_FROM</type>
<position>652,-30</position>
<input>
<ID>IN_0</ID>631 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_ES</lparam></gate>
<gate>
<ID>767</ID>
<type>DA_FROM</type>
<position>652,-33</position>
<input>
<ID>IN_0</ID>632 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_RAM</lparam></gate>
<gate>
<ID>768</ID>
<type>DE_TO</type>
<position>662,-31</position>
<input>
<ID>IN_0</ID>633 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4_MUX_OUT</lparam></gate>
<gate>
<ID>769</ID>
<type>DA_FROM</type>
<position>652,-27</position>
<input>
<ID>IN_0</ID>634 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>770</ID>
<type>AA_MUX_2x1</type>
<position>657,-40</position>
<input>
<ID>IN_0</ID>636 </input>
<input>
<ID>IN_1</ID>635 </input>
<output>
<ID>OUT</ID>637 </output>
<input>
<ID>SEL_0</ID>638 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>771</ID>
<type>DA_FROM</type>
<position>652,-39</position>
<input>
<ID>IN_0</ID>635 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5_ES</lparam></gate>
<wire>
<ID>615</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>654,7,655,7</points>
<connection>
<GID>741</GID>
<name>IN_1</name></connection>
<connection>
<GID>743</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>654,4,654,5</points>
<connection>
<GID>745</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,5,655,5</points>
<connection>
<GID>741</GID>
<name>IN_0</name></connection>
<intersection>654 0</intersection></hsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>659,6,660,6</points>
<connection>
<GID>741</GID>
<name>OUT</name></connection>
<connection>
<GID>747</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>657,8.5,657,10</points>
<connection>
<GID>741</GID>
<name>SEL_0</name></connection>
<intersection>10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,10,657,10</points>
<connection>
<GID>749</GID>
<name>IN_0</name></connection>
<intersection>657 0</intersection></hsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>654,-3,655,-3</points>
<connection>
<GID>750</GID>
<name>IN_1</name></connection>
<connection>
<GID>751</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>654,-6,654,-5</points>
<connection>
<GID>752</GID>
<name>IN_0</name></connection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,-5,655,-5</points>
<connection>
<GID>750</GID>
<name>IN_0</name></connection>
<intersection>654 0</intersection></hsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>659,-4,660,-4</points>
<connection>
<GID>750</GID>
<name>OUT</name></connection>
<connection>
<GID>753</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>657,-1.5,657,0</points>
<connection>
<GID>750</GID>
<name>SEL_0</name></connection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,0,657,0</points>
<connection>
<GID>754</GID>
<name>IN_0</name></connection>
<intersection>657 0</intersection></hsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>654,-12,655,-12</points>
<connection>
<GID>755</GID>
<name>IN_1</name></connection>
<connection>
<GID>756</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>654,-15,654,-14</points>
<connection>
<GID>757</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,-14,655,-14</points>
<connection>
<GID>755</GID>
<name>IN_0</name></connection>
<intersection>654 0</intersection></hsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>659,-13,660,-13</points>
<connection>
<GID>755</GID>
<name>OUT</name></connection>
<connection>
<GID>758</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>657,-10.5,657,-9</points>
<connection>
<GID>755</GID>
<name>SEL_0</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,-9,657,-9</points>
<connection>
<GID>759</GID>
<name>IN_0</name></connection>
<intersection>657 0</intersection></hsegment></shape></wire>
<wire>
<ID>627</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>654,-21,655,-21</points>
<connection>
<GID>760</GID>
<name>IN_1</name></connection>
<connection>
<GID>761</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>628</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>654,-24,654,-23</points>
<connection>
<GID>762</GID>
<name>IN_0</name></connection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,-23,655,-23</points>
<connection>
<GID>760</GID>
<name>IN_0</name></connection>
<intersection>654 0</intersection></hsegment></shape></wire>
<wire>
<ID>629</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>659,-22,660,-22</points>
<connection>
<GID>760</GID>
<name>OUT</name></connection>
<connection>
<GID>763</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>630</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>657,-19.5,657,-18</points>
<connection>
<GID>760</GID>
<name>SEL_0</name></connection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,-18,657,-18</points>
<connection>
<GID>764</GID>
<name>IN_0</name></connection>
<intersection>657 0</intersection></hsegment></shape></wire>
<wire>
<ID>631</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>654,-30,655,-30</points>
<connection>
<GID>765</GID>
<name>IN_1</name></connection>
<connection>
<GID>766</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>632</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>654,-33,654,-32</points>
<connection>
<GID>767</GID>
<name>IN_0</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,-32,655,-32</points>
<connection>
<GID>765</GID>
<name>IN_0</name></connection>
<intersection>654 0</intersection></hsegment></shape></wire>
<wire>
<ID>633</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>659,-31,660,-31</points>
<connection>
<GID>765</GID>
<name>OUT</name></connection>
<connection>
<GID>768</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>634</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>657,-28.5,657,-27</points>
<connection>
<GID>765</GID>
<name>SEL_0</name></connection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,-27,657,-27</points>
<connection>
<GID>769</GID>
<name>IN_0</name></connection>
<intersection>657 0</intersection></hsegment></shape></wire>
<wire>
<ID>635</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>654,-39,655,-39</points>
<connection>
<GID>770</GID>
<name>IN_1</name></connection>
<connection>
<GID>771</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>636</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>654,-42,654,-41</points>
<connection>
<GID>772</GID>
<name>IN_0</name></connection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,-41,655,-41</points>
<connection>
<GID>770</GID>
<name>IN_0</name></connection>
<intersection>654 0</intersection></hsegment></shape></wire>
<wire>
<ID>637</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>659,-40,660,-40</points>
<connection>
<GID>770</GID>
<name>OUT</name></connection>
<connection>
<GID>773</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>638</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>657,-37.5,657,-36</points>
<connection>
<GID>770</GID>
<name>SEL_0</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,-36,657,-36</points>
<connection>
<GID>774</GID>
<name>IN_0</name></connection>
<intersection>657 0</intersection></hsegment></shape></wire>
<wire>
<ID>639</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>654,-48,655,-48</points>
<connection>
<GID>775</GID>
<name>IN_1</name></connection>
<connection>
<GID>776</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>654,-51,654,-50</points>
<connection>
<GID>777</GID>
<name>IN_0</name></connection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,-50,655,-50</points>
<connection>
<GID>775</GID>
<name>IN_0</name></connection>
<intersection>654 0</intersection></hsegment></shape></wire>
<wire>
<ID>641</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>659,-49,660,-49</points>
<connection>
<GID>775</GID>
<name>OUT</name></connection>
<connection>
<GID>778</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>642</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>657,-46.5,657,-45</points>
<connection>
<GID>775</GID>
<name>SEL_0</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,-45,657,-45</points>
<connection>
<GID>779</GID>
<name>IN_0</name></connection>
<intersection>657 0</intersection></hsegment></shape></wire>
<wire>
<ID>643</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>654,-57,655,-57</points>
<connection>
<GID>780</GID>
<name>IN_1</name></connection>
<connection>
<GID>781</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>644</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>654,-60,654,-59</points>
<connection>
<GID>782</GID>
<name>IN_0</name></connection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,-59,655,-59</points>
<connection>
<GID>780</GID>
<name>IN_0</name></connection>
<intersection>654 0</intersection></hsegment></shape></wire>
<wire>
<ID>645</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>659,-58,660,-58</points>
<connection>
<GID>780</GID>
<name>OUT</name></connection>
<connection>
<GID>783</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>646</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>657,-55.5,657,-54</points>
<connection>
<GID>780</GID>
<name>SEL_0</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,-54,657,-54</points>
<connection>
<GID>784</GID>
<name>IN_0</name></connection>
<intersection>657 0</intersection></hsegment></shape></wire>
<wire>
<ID>647</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>714,6.5,715,6.5</points>
<connection>
<GID>785</GID>
<name>IN_1</name></connection>
<connection>
<GID>786</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>648</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>714,3.5,714,4.5</points>
<connection>
<GID>787</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,4.5,715,4.5</points>
<connection>
<GID>785</GID>
<name>IN_0</name></connection>
<intersection>714 0</intersection></hsegment></shape></wire>
<wire>
<ID>649</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>719,5.5,720,5.5</points>
<connection>
<GID>785</GID>
<name>OUT</name></connection>
<connection>
<GID>788</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>650</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>717,8,717,9.5</points>
<connection>
<GID>785</GID>
<name>SEL_0</name></connection>
<intersection>9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,9.5,717,9.5</points>
<connection>
<GID>789</GID>
<name>IN_0</name></connection>
<intersection>717 0</intersection></hsegment></shape></wire>
<wire>
<ID>651</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>714,-2.5,715,-2.5</points>
<connection>
<GID>790</GID>
<name>IN_1</name></connection>
<connection>
<GID>791</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>652</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>714,-5.5,714,-4.5</points>
<connection>
<GID>792</GID>
<name>IN_0</name></connection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,-4.5,715,-4.5</points>
<connection>
<GID>790</GID>
<name>IN_0</name></connection>
<intersection>714 0</intersection></hsegment></shape></wire>
<wire>
<ID>653</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>719,-3.5,720,-3.5</points>
<connection>
<GID>790</GID>
<name>OUT</name></connection>
<connection>
<GID>793</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>654</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>717,-1,717,0.5</points>
<connection>
<GID>790</GID>
<name>SEL_0</name></connection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,0.5,717,0.5</points>
<connection>
<GID>794</GID>
<name>IN_0</name></connection>
<intersection>717 0</intersection></hsegment></shape></wire>
<wire>
<ID>655</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>714,-11.5,715,-11.5</points>
<connection>
<GID>795</GID>
<name>IN_1</name></connection>
<connection>
<GID>796</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>656</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>714,-14.5,714,-13.5</points>
<connection>
<GID>797</GID>
<name>IN_0</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,-13.5,715,-13.5</points>
<connection>
<GID>795</GID>
<name>IN_0</name></connection>
<intersection>714 0</intersection></hsegment></shape></wire>
<wire>
<ID>657</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>719,-12.5,720,-12.5</points>
<connection>
<GID>795</GID>
<name>OUT</name></connection>
<connection>
<GID>798</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>658</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>717,-10,717,-8.5</points>
<connection>
<GID>795</GID>
<name>SEL_0</name></connection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,-8.5,717,-8.5</points>
<connection>
<GID>799</GID>
<name>IN_0</name></connection>
<intersection>717 0</intersection></hsegment></shape></wire>
<wire>
<ID>659</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>714,-20.5,715,-20.5</points>
<connection>
<GID>800</GID>
<name>IN_1</name></connection>
<connection>
<GID>801</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>660</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>714,-23.5,714,-22.5</points>
<connection>
<GID>802</GID>
<name>IN_0</name></connection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,-22.5,715,-22.5</points>
<connection>
<GID>800</GID>
<name>IN_0</name></connection>
<intersection>714 0</intersection></hsegment></shape></wire>
<wire>
<ID>661</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>719,-21.5,720,-21.5</points>
<connection>
<GID>800</GID>
<name>OUT</name></connection>
<connection>
<GID>803</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>662</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>717,-19,717,-17.5</points>
<connection>
<GID>800</GID>
<name>SEL_0</name></connection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,-17.5,717,-17.5</points>
<connection>
<GID>804</GID>
<name>IN_0</name></connection>
<intersection>717 0</intersection></hsegment></shape></wire>
<wire>
<ID>663</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>714,-29.5,715,-29.5</points>
<connection>
<GID>805</GID>
<name>IN_1</name></connection>
<connection>
<GID>806</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>664</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>714,-32.5,714,-31.5</points>
<connection>
<GID>807</GID>
<name>IN_0</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,-31.5,715,-31.5</points>
<connection>
<GID>805</GID>
<name>IN_0</name></connection>
<intersection>714 0</intersection></hsegment></shape></wire>
<wire>
<ID>665</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>719,-30.5,720,-30.5</points>
<connection>
<GID>805</GID>
<name>OUT</name></connection>
<connection>
<GID>808</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>717,-28,717,-26.5</points>
<connection>
<GID>805</GID>
<name>SEL_0</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,-26.5,717,-26.5</points>
<connection>
<GID>809</GID>
<name>IN_0</name></connection>
<intersection>717 0</intersection></hsegment></shape></wire>
<wire>
<ID>667</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>714,-38.5,715,-38.5</points>
<connection>
<GID>810</GID>
<name>IN_1</name></connection>
<connection>
<GID>811</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>668</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>714,-41.5,714,-40.5</points>
<connection>
<GID>812</GID>
<name>IN_0</name></connection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,-40.5,715,-40.5</points>
<connection>
<GID>810</GID>
<name>IN_0</name></connection>
<intersection>714 0</intersection></hsegment></shape></wire>
<wire>
<ID>669</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>719,-39.5,720,-39.5</points>
<connection>
<GID>810</GID>
<name>OUT</name></connection>
<connection>
<GID>813</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>670</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>717,-37,717,-35.5</points>
<connection>
<GID>810</GID>
<name>SEL_0</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,-35.5,717,-35.5</points>
<connection>
<GID>814</GID>
<name>IN_0</name></connection>
<intersection>717 0</intersection></hsegment></shape></wire>
<wire>
<ID>671</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>714,-47.5,715,-47.5</points>
<connection>
<GID>815</GID>
<name>IN_1</name></connection>
<connection>
<GID>816</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>672</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>714,-50.5,714,-49.5</points>
<connection>
<GID>817</GID>
<name>IN_0</name></connection>
<intersection>-49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,-49.5,715,-49.5</points>
<connection>
<GID>815</GID>
<name>IN_0</name></connection>
<intersection>714 0</intersection></hsegment></shape></wire>
<wire>
<ID>673</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>719,-48.5,720,-48.5</points>
<connection>
<GID>815</GID>
<name>OUT</name></connection>
<connection>
<GID>818</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>674</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>717,-46,717,-44.5</points>
<connection>
<GID>815</GID>
<name>SEL_0</name></connection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,-44.5,717,-44.5</points>
<connection>
<GID>819</GID>
<name>IN_0</name></connection>
<intersection>717 0</intersection></hsegment></shape></wire>
<wire>
<ID>675</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>714,-56.5,715,-56.5</points>
<connection>
<GID>820</GID>
<name>IN_1</name></connection>
<connection>
<GID>821</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>676</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>714,-59.5,714,-58.5</points>
<connection>
<GID>822</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,-58.5,715,-58.5</points>
<connection>
<GID>820</GID>
<name>IN_0</name></connection>
<intersection>714 0</intersection></hsegment></shape></wire>
<wire>
<ID>677</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>719,-57.5,720,-57.5</points>
<connection>
<GID>820</GID>
<name>OUT</name></connection>
<connection>
<GID>823</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>678</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>717,-55,717,-53.5</points>
<connection>
<GID>820</GID>
<name>SEL_0</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,-53.5,717,-53.5</points>
<connection>
<GID>824</GID>
<name>IN_0</name></connection>
<intersection>717 0</intersection></hsegment></shape></wire></page 6>
<page 7>
<PageViewport>589.739,40.3387,799.353,-67.7688</PageViewport>
<gate>
<ID>969</ID>
<type>AE_OR4</type>
<position>643,-8</position>
<input>
<ID>IN_0</ID>811 </input>
<input>
<ID>IN_1</ID>813 </input>
<input>
<ID>IN_2</ID>814 </input>
<input>
<ID>IN_3</ID>815 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>970</ID>
<type>DA_FROM</type>
<position>626,-13</position>
<input>
<ID>IN_0</ID>815 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15_IR</lparam></gate>
<gate>
<ID>1017</ID>
<type>AA_LABEL</type>
<position>672,38.5</position>
<gparam>LABEL_TEXT Decodificador de Instrucoes</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>828</ID>
<type>AA_AND3</type>
<position>635.5,25.5</position>
<input>
<ID>IN_0</ID>686 </input>
<input>
<ID>IN_1</ID>687 </input>
<input>
<ID>IN_2</ID>688 </input>
<output>
<ID>OUT</ID>1037 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>829</ID>
<type>DA_FROM</type>
<position>626,28.5</position>
<input>
<ID>IN_0</ID>686 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D15_IR</lparam></gate>
<gate>
<ID>830</ID>
<type>DA_FROM</type>
<position>626,25.5</position>
<input>
<ID>IN_0</ID>687 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_IR</lparam></gate>
<gate>
<ID>831</ID>
<type>DA_FROM</type>
<position>626,22</position>
<input>
<ID>IN_0</ID>688 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_IR</lparam></gate>
<gate>
<ID>836</ID>
<type>DA_FROM</type>
<position>692,5.5</position>
<input>
<ID>IN_0</ID>1033 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D15_IR</lparam></gate>
<gate>
<ID>837</ID>
<type>DA_FROM</type>
<position>692,2</position>
<input>
<ID>IN_0</ID>1034 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D14_IR</lparam></gate>
<gate>
<ID>838</ID>
<type>DA_FROM</type>
<position>692,-2</position>
<input>
<ID>IN_0</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D13_IR</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_LABEL</type>
<position>663.5,55</position>
<gparam>LABEL_TEXT Prof.  Angelo Zanini / Nuncio Perrella</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>270</ID>
<type>AA_LABEL</type>
<position>661.5,64.5</position>
<gparam>LABEL_TEXT PROCESSADOR BIP IMT - MAUA 2022</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_INVERTER</type>
<position>643,2</position>
<input>
<ID>IN_0</ID>56 </input>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>892</ID>
<type>AA_AND4</type>
<position>701.5,13.5</position>
<input>
<ID>IN_0</ID>739 </input>
<input>
<ID>IN_1</ID>740 </input>
<input>
<ID>IN_2</ID>741 </input>
<input>
<ID>IN_3</ID>742 </input>
<output>
<ID>OUT</ID>1076 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>894</ID>
<type>DA_FROM</type>
<position>692,18.5</position>
<input>
<ID>IN_0</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D15_IR</lparam></gate>
<gate>
<ID>895</ID>
<type>DA_FROM</type>
<position>692,15</position>
<input>
<ID>IN_0</ID>740 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D14_IR</lparam></gate>
<gate>
<ID>896</ID>
<type>DA_FROM</type>
<position>692,12</position>
<input>
<ID>IN_0</ID>741 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_IR</lparam></gate>
<gate>
<ID>897</ID>
<type>DA_FROM</type>
<position>692,9</position>
<input>
<ID>IN_0</ID>742 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_IR</lparam></gate>
<gate>
<ID>905</ID>
<type>DE_TO</type>
<position>655,25.5</position>
<input>
<ID>IN_0</ID>1037 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelUlaSrc</lparam></gate>
<gate>
<ID>1299</ID>
<type>AA_AND2</type>
<position>702,4</position>
<input>
<ID>IN_0</ID>1033 </input>
<input>
<ID>IN_1</ID>1034 </input>
<output>
<ID>OUT</ID>1031 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1301</ID>
<type>AA_AND2</type>
<position>702,-3</position>
<input>
<ID>IN_0</ID>1036 </input>
<input>
<ID>IN_1</ID>1035 </input>
<output>
<ID>OUT</ID>1032 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1303</ID>
<type>AE_OR2</type>
<position>710,1</position>
<input>
<ID>IN_0</ID>1031 </input>
<input>
<ID>IN_1</ID>1032 </input>
<output>
<ID>OUT</ID>1059 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>917</ID>
<type>DE_TO</type>
<position>719,1</position>
<input>
<ID>IN_0</ID>1059 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP_ULA</lparam></gate>
<gate>
<ID>1304</ID>
<type>DA_FROM</type>
<position>692,-5.5</position>
<input>
<ID>IN_0</ID>1035 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D15_IR</lparam></gate>
<gate>
<ID>918</ID>
<type>AA_AND3</type>
<position>635,14.5</position>
<input>
<ID>IN_0</ID>721 </input>
<input>
<ID>IN_1</ID>722 </input>
<input>
<ID>IN_2</ID>723 </input>
<output>
<ID>OUT</ID>725 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>919</ID>
<type>DA_FROM</type>
<position>626,18</position>
<input>
<ID>IN_0</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D15_IR</lparam></gate>
<gate>
<ID>920</ID>
<type>DA_FROM</type>
<position>626,14.5</position>
<input>
<ID>IN_0</ID>722 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D14_IR</lparam></gate>
<gate>
<ID>921</ID>
<type>DA_FROM</type>
<position>626,10.5</position>
<input>
<ID>IN_0</ID>723 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D13_IR</lparam></gate>
<gate>
<ID>922</ID>
<type>DE_TO</type>
<position>655,13.5</position>
<input>
<ID>IN_0</ID>726 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WR_RAM</lparam></gate>
<gate>
<ID>924</ID>
<type>AA_AND2</type>
<position>643.5,13.5</position>
<input>
<ID>IN_0</ID>725 </input>
<input>
<ID>IN_1</ID>727 </input>
<output>
<ID>OUT</ID>726 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>925</ID>
<type>DA_FROM</type>
<position>626,7</position>
<input>
<ID>IN_0</ID>727 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_IR</lparam></gate>
<gate>
<ID>926</ID>
<type>DA_FROM</type>
<position>626,2</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>929</ID>
<type>DE_TO</type>
<position>665,-9</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WR_PC</lparam></gate>
<gate>
<ID>931</ID>
<type>DE_TO</type>
<position>655,2</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WR_IR</lparam></gate>
<gate>
<ID>937</ID>
<type>DA_FROM</type>
<position>626,-4</position>
<input>
<ID>IN_0</ID>811 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_IR</lparam></gate>
<gate>
<ID>938</ID>
<type>DE_TO</type>
<position>655.5,-22</position>
<input>
<ID>IN_0</ID>1072 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WR_ACC</lparam></gate>
<gate>
<ID>941</ID>
<type>DA_FROM</type>
<position>626,-7</position>
<input>
<ID>IN_0</ID>813 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12_IR</lparam></gate>
<gate>
<ID>1328</ID>
<type>DA_FROM</type>
<position>626,-17</position>
<input>
<ID>IN_0</ID>1062 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D15_IR</lparam></gate>
<gate>
<ID>1329</ID>
<type>DA_FROM</type>
<position>626,-20.5</position>
<input>
<ID>IN_0</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_IR</lparam></gate>
<gate>
<ID>943</ID>
<type>DA_FROM</type>
<position>626,-10</position>
<input>
<ID>IN_0</ID>814 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_IR</lparam></gate>
<gate>
<ID>1330</ID>
<type>DA_FROM</type>
<position>626,-24.5</position>
<input>
<ID>IN_0</ID>1065 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13_IR</lparam></gate>
<gate>
<ID>1331</ID>
<type>AA_AND2</type>
<position>637.5,-18.5</position>
<input>
<ID>IN_0</ID>1062 </input>
<input>
<ID>IN_1</ID>1063 </input>
<output>
<ID>OUT</ID>1060 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1332</ID>
<type>AA_AND2</type>
<position>637.5,-26.5</position>
<input>
<ID>IN_0</ID>1065 </input>
<input>
<ID>IN_1</ID>1064 </input>
<output>
<ID>OUT</ID>1061 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>946</ID>
<type>DE_TO</type>
<position>717,13.5</position>
<input>
<ID>IN_0</ID>1076 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_0</lparam></gate>
<gate>
<ID>1333</ID>
<type>AE_OR2</type>
<position>647.5,-22</position>
<input>
<ID>IN_0</ID>1060 </input>
<input>
<ID>IN_1</ID>1061 </input>
<output>
<ID>OUT</ID>1072 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1334</ID>
<type>DA_FROM</type>
<position>625.5,-28</position>
<input>
<ID>IN_0</ID>1064 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D15_IR</lparam></gate>
<gate>
<ID>948</ID>
<type>DA_FROM</type>
<position>692,26</position>
<input>
<ID>IN_0</ID>1073 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D15_IR</lparam></gate>
<gate>
<ID>949</ID>
<type>DA_FROM</type>
<position>692,22.5</position>
<input>
<ID>IN_0</ID>1074 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14_IR</lparam></gate>
<gate>
<ID>1336</ID>
<type>AA_AND2</type>
<position>703.5,24.5</position>
<input>
<ID>IN_0</ID>1073 </input>
<input>
<ID>IN_1</ID>1074 </input>
<output>
<ID>OUT</ID>1075 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>951</ID>
<type>DE_TO</type>
<position>717,24.5</position>
<input>
<ID>IN_0</ID>1075 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SelAccSrc_1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>655,-9,655,-8</points>
<intersection>-9 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>655,-9,663,-9</points>
<connection>
<GID>929</GID>
<name>IN_0</name></connection>
<intersection>655 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>647,-8,655,-8</points>
<connection>
<GID>969</GID>
<name>OUT</name></connection>
<intersection>655 0</intersection></hsegment></shape></wire>
<wire>
<ID>811</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>631,-5,631,-4</points>
<intersection>-5 1</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>631,-5,640,-5</points>
<connection>
<GID>969</GID>
<name>IN_0</name></connection>
<intersection>631 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>628,-4,631,-4</points>
<connection>
<GID>937</GID>
<name>IN_0</name></connection>
<intersection>631 0</intersection></hsegment></shape></wire>
<wire>
<ID>813</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>628,-7,640,-7</points>
<connection>
<GID>941</GID>
<name>IN_0</name></connection>
<connection>
<GID>969</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>814</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>632.5,-10,632.5,-9</points>
<intersection>-10 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>632.5,-9,640,-9</points>
<connection>
<GID>969</GID>
<name>IN_2</name></connection>
<intersection>632.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>628,-10,632.5,-10</points>
<connection>
<GID>943</GID>
<name>IN_0</name></connection>
<intersection>632.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>815</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>634,-13,634,-11</points>
<intersection>-13 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>634,-11,640,-11</points>
<connection>
<GID>969</GID>
<name>IN_3</name></connection>
<intersection>634 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>628,-13,634,-13</points>
<connection>
<GID>970</GID>
<name>IN_0</name></connection>
<intersection>634 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>628,2,640,2</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<connection>
<GID>926</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1031</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>706,2,707,2</points>
<connection>
<GID>1303</GID>
<name>IN_0</name></connection>
<intersection>706 1</intersection></hsegment>
<vsegment>
<ID>1</ID>
<points>706,2,706,4</points>
<intersection>2 0</intersection>
<intersection>4 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>705,4,706,4</points>
<connection>
<GID>1299</GID>
<name>OUT</name></connection>
<intersection>706 1</intersection></hsegment></shape></wire>
<wire>
<ID>1032</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>706,-3,706,0</points>
<intersection>-3 1</intersection>
<intersection>0 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>705,-3,706,-3</points>
<connection>
<GID>1301</GID>
<name>OUT</name></connection>
<intersection>706 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>706,0,707,0</points>
<connection>
<GID>1303</GID>
<name>IN_1</name></connection>
<intersection>706 0</intersection></hsegment></shape></wire>
<wire>
<ID>1033</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>697,5,697,5.5</points>
<intersection>5 1</intersection>
<intersection>5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>697,5,699,5</points>
<connection>
<GID>1299</GID>
<name>IN_0</name></connection>
<intersection>697 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>694,5.5,697,5.5</points>
<connection>
<GID>836</GID>
<name>IN_0</name></connection>
<intersection>697 0</intersection></hsegment></shape></wire>
<wire>
<ID>1034</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>697,2,697,3</points>
<intersection>2 2</intersection>
<intersection>3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>697,3,699,3</points>
<connection>
<GID>1299</GID>
<name>IN_1</name></connection>
<intersection>697 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>694,2,697,2</points>
<connection>
<GID>837</GID>
<name>IN_0</name></connection>
<intersection>697 0</intersection></hsegment></shape></wire>
<wire>
<ID>1035</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>697,-5.5,697,-4</points>
<intersection>-5.5 2</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>697,-4,699,-4</points>
<connection>
<GID>1301</GID>
<name>IN_1</name></connection>
<intersection>697 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>694,-5.5,697,-5.5</points>
<connection>
<GID>1304</GID>
<name>IN_0</name></connection>
<intersection>697 0</intersection></hsegment></shape></wire>
<wire>
<ID>1036</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>694,-2,699,-2</points>
<connection>
<GID>838</GID>
<name>IN_0</name></connection>
<connection>
<GID>1301</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1037</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>638.5,25.5,653,25.5</points>
<connection>
<GID>828</GID>
<name>OUT</name></connection>
<connection>
<GID>905</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>646,2,653,2</points>
<connection>
<GID>931</GID>
<name>IN_0</name></connection>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1059</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>713,1,717,1</points>
<connection>
<GID>1303</GID>
<name>OUT</name></connection>
<connection>
<GID>917</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1060</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>642.5,-21,644.5,-21</points>
<connection>
<GID>1333</GID>
<name>IN_0</name></connection>
<intersection>642.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>642.5,-21,642.5,-18.5</points>
<intersection>-21 1</intersection>
<intersection>-18.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>640.5,-18.5,642.5,-18.5</points>
<connection>
<GID>1331</GID>
<name>OUT</name></connection>
<intersection>642.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1061</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>642.5,-26.5,642.5,-23</points>
<intersection>-26.5 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640.5,-26.5,642.5,-26.5</points>
<connection>
<GID>1332</GID>
<name>OUT</name></connection>
<intersection>642.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>642.5,-23,644.5,-23</points>
<connection>
<GID>1333</GID>
<name>IN_1</name></connection>
<intersection>642.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1062</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>631,-17.5,631,-17</points>
<intersection>-17.5 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>631,-17.5,634.5,-17.5</points>
<connection>
<GID>1331</GID>
<name>IN_0</name></connection>
<intersection>631 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>628,-17,631,-17</points>
<connection>
<GID>1328</GID>
<name>IN_0</name></connection>
<intersection>631 0</intersection></hsegment></shape></wire>
<wire>
<ID>1063</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>631,-20.5,631,-19.5</points>
<intersection>-20.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>631,-19.5,634.5,-19.5</points>
<connection>
<GID>1331</GID>
<name>IN_1</name></connection>
<intersection>631 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>628,-20.5,631,-20.5</points>
<connection>
<GID>1329</GID>
<name>IN_0</name></connection>
<intersection>631 0</intersection></hsegment></shape></wire>
<wire>
<ID>1064</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>631,-28,631,-27.5</points>
<intersection>-28 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>631,-27.5,634.5,-27.5</points>
<connection>
<GID>1332</GID>
<name>IN_1</name></connection>
<intersection>631 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>627.5,-28,631,-28</points>
<connection>
<GID>1334</GID>
<name>IN_0</name></connection>
<intersection>631 0</intersection></hsegment></shape></wire>
<wire>
<ID>1065</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>631,-25.5,631,-24.5</points>
<intersection>-25.5 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>631,-25.5,634.5,-25.5</points>
<connection>
<GID>1332</GID>
<name>IN_0</name></connection>
<intersection>631 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>628,-24.5,631,-24.5</points>
<connection>
<GID>1330</GID>
<name>IN_0</name></connection>
<intersection>631 0</intersection></hsegment></shape></wire>
<wire>
<ID>1072</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>650.5,-22,653.5,-22</points>
<connection>
<GID>1333</GID>
<name>OUT</name></connection>
<connection>
<GID>938</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>686</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>628,28.5,632,28.5</points>
<connection>
<GID>829</GID>
<name>IN_0</name></connection>
<intersection>632 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>632,27.5,632,28.5</points>
<intersection>27.5 5</intersection>
<intersection>28.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>632,27.5,632.5,27.5</points>
<connection>
<GID>828</GID>
<name>IN_0</name></connection>
<intersection>632 3</intersection></hsegment></shape></wire>
<wire>
<ID>1073</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>697,25.5,697,26</points>
<intersection>25.5 1</intersection>
<intersection>26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>697,25.5,700.5,25.5</points>
<connection>
<GID>1336</GID>
<name>IN_0</name></connection>
<intersection>697 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>694,26,697,26</points>
<connection>
<GID>948</GID>
<name>IN_0</name></connection>
<intersection>697 0</intersection></hsegment></shape></wire>
<wire>
<ID>687</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>628,25.5,632.5,25.5</points>
<connection>
<GID>828</GID>
<name>IN_1</name></connection>
<connection>
<GID>830</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1074</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>697,22.5,697,23.5</points>
<intersection>22.5 2</intersection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>697,23.5,700.5,23.5</points>
<connection>
<GID>1336</GID>
<name>IN_1</name></connection>
<intersection>697 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>694,22.5,697,22.5</points>
<connection>
<GID>949</GID>
<name>IN_0</name></connection>
<intersection>697 0</intersection></hsegment></shape></wire>
<wire>
<ID>688</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>632,22,632,23.5</points>
<intersection>22 2</intersection>
<intersection>23.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>628,22,632,22</points>
<connection>
<GID>831</GID>
<name>IN_0</name></connection>
<intersection>632 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>632,23.5,632.5,23.5</points>
<connection>
<GID>828</GID>
<name>IN_2</name></connection>
<intersection>632 0</intersection></hsegment></shape></wire>
<wire>
<ID>1075</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>706.5,24.5,715,24.5</points>
<connection>
<GID>1336</GID>
<name>OUT</name></connection>
<connection>
<GID>951</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1076</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>704.5,13.5,715,13.5</points>
<connection>
<GID>892</GID>
<name>OUT</name></connection>
<connection>
<GID>946</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>721</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>628,18,629,18</points>
<connection>
<GID>919</GID>
<name>IN_0</name></connection>
<intersection>629 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>629,16.5,629,18</points>
<intersection>16.5 4</intersection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>629,16.5,632,16.5</points>
<connection>
<GID>918</GID>
<name>IN_0</name></connection>
<intersection>629 3</intersection></hsegment></shape></wire>
<wire>
<ID>722</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>628,14.5,632,14.5</points>
<connection>
<GID>920</GID>
<name>IN_0</name></connection>
<connection>
<GID>918</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>723</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>629,10.5,629,12.5</points>
<intersection>10.5 2</intersection>
<intersection>12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>629,12.5,632,12.5</points>
<connection>
<GID>918</GID>
<name>IN_2</name></connection>
<intersection>629 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>628,10.5,629,10.5</points>
<connection>
<GID>921</GID>
<name>IN_0</name></connection>
<intersection>629 0</intersection></hsegment></shape></wire>
<wire>
<ID>725</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>638,14.5,640.5,14.5</points>
<connection>
<GID>924</GID>
<name>IN_0</name></connection>
<connection>
<GID>918</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>726</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>646.5,13.5,653,13.5</points>
<connection>
<GID>924</GID>
<name>OUT</name></connection>
<connection>
<GID>922</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>727</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>638,7,638,12.5</points>
<intersection>7 2</intersection>
<intersection>12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>638,12.5,640.5,12.5</points>
<connection>
<GID>924</GID>
<name>IN_1</name></connection>
<intersection>638 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>628,7,638,7</points>
<connection>
<GID>925</GID>
<name>IN_0</name></connection>
<intersection>638 0</intersection></hsegment></shape></wire>
<wire>
<ID>739</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>694,18.5,697,18.5</points>
<connection>
<GID>894</GID>
<name>IN_0</name></connection>
<intersection>697 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>697,16.5,697,18.5</points>
<intersection>16.5 3</intersection>
<intersection>18.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>697,16.5,698.5,16.5</points>
<connection>
<GID>892</GID>
<name>IN_0</name></connection>
<intersection>697 2</intersection></hsegment></shape></wire>
<wire>
<ID>740</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>696,14.5,696,15</points>
<intersection>14.5 1</intersection>
<intersection>15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>696,14.5,698.5,14.5</points>
<connection>
<GID>892</GID>
<name>IN_1</name></connection>
<intersection>696 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>694,15,696,15</points>
<connection>
<GID>895</GID>
<name>IN_0</name></connection>
<intersection>696 0</intersection></hsegment></shape></wire>
<wire>
<ID>741</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>696,12,696,12.5</points>
<intersection>12 2</intersection>
<intersection>12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>696,12.5,698.5,12.5</points>
<connection>
<GID>892</GID>
<name>IN_2</name></connection>
<intersection>696 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>694,12,696,12</points>
<connection>
<GID>896</GID>
<name>IN_0</name></connection>
<intersection>696 0</intersection></hsegment></shape></wire>
<wire>
<ID>742</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>697.5,9,697.5,10.5</points>
<intersection>9 2</intersection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>697.5,10.5,698.5,10.5</points>
<connection>
<GID>892</GID>
<name>IN_3</name></connection>
<intersection>697.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>694,9,697.5,9</points>
<connection>
<GID>897</GID>
<name>IN_0</name></connection>
<intersection>697.5 0</intersection></hsegment></shape></wire></page 7>
<page 8>
<PageViewport>763.89,665.28,1080.34,502.074</PageViewport>
<gate>
<ID>825</ID>
<type>DA_FROM</type>
<position>893,570.5</position>
<input>
<ID>IN_0</ID>194 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D8_ACC_OUT</lparam></gate>
<gate>
<ID>827</ID>
<type>DE_TO</type>
<position>914,552.5</position>
<input>
<ID>IN_0</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLOCK</lparam></gate>
<gate>
<ID>832</ID>
<type>AA_AND2</type>
<position>898,548.5</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>833</ID>
<type>AE_OR2</type>
<position>905,552.5</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>834</ID>
<type>AA_LABEL</type>
<position>846,554</position>
<gparam>LABEL_TEXT STEP</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>835</ID>
<type>AA_TOGGLE</type>
<position>854,553.5</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>839</ID>
<type>AA_LABEL</type>
<position>846,549.5</position>
<gparam>LABEL_TEXT HALT</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>454</ID>
<type>DA_FROM</type>
<position>914,564.5</position>
<input>
<ID>IN_0</ID>188 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D2_ACC_OUT</lparam></gate>
<gate>
<ID>840</ID>
<type>AA_TOGGLE</type>
<position>853.5,549</position>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>841</ID>
<type>DA_FROM</type>
<position>869,569.5</position>
<input>
<ID>IN_0</ID>212 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PCA0</lparam></gate>
<gate>
<ID>842</ID>
<type>DA_FROM</type>
<position>869,566.5</position>
<input>
<ID>IN_0</ID>217 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PCA1</lparam></gate>
<gate>
<ID>457</ID>
<type>DA_FROM</type>
<position>914,567.5</position>
<input>
<ID>IN_0</ID>187 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D1_ACC_OUT</lparam></gate>
<gate>
<ID>843</ID>
<type>DA_FROM</type>
<position>869,563.5</position>
<input>
<ID>IN_0</ID>220 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PCA2</lparam></gate>
<gate>
<ID>844</ID>
<type>DA_FROM</type>
<position>869,560.5</position>
<input>
<ID>IN_0</ID>221 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PCA3</lparam></gate>
<gate>
<ID>845</ID>
<type>DA_FROM</type>
<position>869,595.5</position>
<input>
<ID>IN_0</ID>254 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PCA4</lparam></gate>
<gate>
<ID>460</ID>
<type>DA_FROM</type>
<position>914,570.5</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D0_ACC_OUT</lparam></gate>
<gate>
<ID>846</ID>
<type>DA_FROM</type>
<position>869,592.5</position>
<input>
<ID>IN_0</ID>250 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PCA5</lparam></gate>
<gate>
<ID>268</ID>
<type>DA_FROM</type>
<position>830.5,561.5</position>
<input>
<ID>IN_0</ID>689 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D15_IR</lparam></gate>
<gate>
<ID>847</ID>
<type>AA_LABEL</type>
<position>847,545.5</position>
<gparam>LABEL_TEXT RESET</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>848</ID>
<type>DA_FROM</type>
<position>869,589.5</position>
<input>
<ID>IN_0</ID>246 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PCA6</lparam></gate>
<gate>
<ID>271</ID>
<type>AA_LABEL</type>
<position>835,604</position>
<gparam>LABEL_TEXT Instrucao</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>850</ID>
<type>DA_FROM</type>
<position>869,586.5</position>
<input>
<ID>IN_0</ID>245 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PCA7</lparam></gate>
<gate>
<ID>273</ID>
<type>AA_LABEL</type>
<position>908,603.5</position>
<gparam>LABEL_TEXT Acumulador</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>857</ID>
<type>BB_CLOCK</type>
<position>886.5,546</position>
<output>
<ID>CLK</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 10</lparam></gate>
<gate>
<ID>859</ID>
<type>DA_FROM</type>
<position>853.5,569.5</position>
<input>
<ID>IN_0</ID>679 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PCA8</lparam></gate>
<gate>
<ID>281</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>920.5,578</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>187 </input>
<input>
<ID>IN_2</ID>188 </input>
<input>
<ID>IN_3</ID>189 </input>
<input>
<ID>IN_4</ID>69 </input>
<input>
<ID>IN_5</ID>68 </input>
<input>
<ID>IN_6</ID>67 </input>
<input>
<ID>IN_7</ID>66 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 83</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>864</ID>
<type>DA_FROM</type>
<position>853.5,566.5</position>
<input>
<ID>IN_0</ID>680 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PCA9</lparam></gate>
<gate>
<ID>865</ID>
<type>DA_FROM</type>
<position>853.5,563.5</position>
<input>
<ID>IN_0</ID>681 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PCA10</lparam></gate>
<gate>
<ID>481</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>899.5,578</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>195 </input>
<input>
<ID>IN_2</ID>196 </input>
<input>
<ID>IN_3</ID>208 </input>
<input>
<ID>IN_4</ID>193 </input>
<input>
<ID>IN_5</ID>192 </input>
<input>
<ID>IN_6</ID>191 </input>
<input>
<ID>IN_7</ID>190 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>867</ID>
<type>DA_FROM</type>
<position>853.5,560.5</position>
<input>
<ID>IN_0</ID>682 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PCA11</lparam></gate>
<gate>
<ID>870</ID>
<type>AA_TOGGLE</type>
<position>854,545.5</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>873</ID>
<type>DE_TO</type>
<position>859.5,545.5</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RESET</lparam></gate>
<gate>
<ID>295</ID>
<type>DA_FROM</type>
<position>914,586.5</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D7_ACC_OUT</lparam></gate>
<gate>
<ID>299</ID>
<type>DA_FROM</type>
<position>914,589.5</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D6_ACC_OUT</lparam></gate>
<gate>
<ID>310</ID>
<type>DA_FROM</type>
<position>914,592.5</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D5_ACC_OUT</lparam></gate>
<gate>
<ID>311</ID>
<type>DA_FROM</type>
<position>914,595.5</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D4_ACC_OUT</lparam></gate>
<gate>
<ID>890</ID>
<type>AA_LABEL</type>
<position>864,603</position>
<gparam>LABEL_TEXT PC </gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>312</ID>
<type>DA_FROM</type>
<position>914,561.5</position>
<input>
<ID>IN_0</ID>189 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D3_ACC_OUT</lparam></gate>
<gate>
<ID>893</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>833.5,578</position>
<input>
<ID>IN_0</ID>683 </input>
<input>
<ID>IN_1</ID>684 </input>
<input>
<ID>IN_2</ID>685 </input>
<input>
<ID>IN_3</ID>689 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>898</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>872,577.5</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>217 </input>
<input>
<ID>IN_2</ID>220 </input>
<input>
<ID>IN_3</ID>221 </input>
<input>
<ID>IN_4</ID>254 </input>
<input>
<ID>IN_5</ID>250 </input>
<input>
<ID>IN_6</ID>246 </input>
<input>
<ID>IN_7</ID>245 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 26</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>899</ID>
<type>DA_FROM</type>
<position>830.5,570.5</position>
<input>
<ID>IN_0</ID>683 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D12_IR</lparam></gate>
<gate>
<ID>900</ID>
<type>DA_FROM</type>
<position>830.5,567.5</position>
<input>
<ID>IN_0</ID>684 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D13_IR</lparam></gate>
<gate>
<ID>901</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>856.5,577.5</position>
<input>
<ID>IN_0</ID>679 </input>
<input>
<ID>IN_1</ID>680 </input>
<input>
<ID>IN_2</ID>681 </input>
<input>
<ID>IN_3</ID>682 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>902</ID>
<type>DA_FROM</type>
<position>830.5,564.5</position>
<input>
<ID>IN_0</ID>685 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D14_IR</lparam></gate>
<gate>
<ID>903</ID>
<type>AA_LABEL</type>
<position>876.5,630.5</position>
<gparam>LABEL_TEXT PROCESSADOR BIP IMT - MAUA 2022</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>904</ID>
<type>AA_LABEL</type>
<position>870,620.5</position>
<gparam>LABEL_TEXT Prof.  Angelo Zanini / Nuncio Perrella</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>736</ID>
<type>DA_FROM</type>
<position>893,586.5</position>
<input>
<ID>IN_0</ID>190 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D15_ACC_OUT</lparam></gate>
<gate>
<ID>738</ID>
<type>DA_FROM</type>
<position>893,589.5</position>
<input>
<ID>IN_0</ID>191 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D14_ACC_OUT</lparam></gate>
<gate>
<ID>740</ID>
<type>DA_FROM</type>
<position>893,592.5</position>
<input>
<ID>IN_0</ID>192 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D13_ACC_OUT</lparam></gate>
<gate>
<ID>742</ID>
<type>DA_FROM</type>
<position>893,595.5</position>
<input>
<ID>IN_0</ID>193 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D12_ACC_OUT</lparam></gate>
<gate>
<ID>744</ID>
<type>DA_FROM</type>
<position>893,561.5</position>
<input>
<ID>IN_0</ID>208 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D11_ACC_OUT</lparam></gate>
<gate>
<ID>746</ID>
<type>DA_FROM</type>
<position>893,564.5</position>
<input>
<ID>IN_0</ID>196 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D10_ACC_OUT</lparam></gate>
<gate>
<ID>748</ID>
<type>DA_FROM</type>
<position>893,567.5</position>
<input>
<ID>IN_0</ID>195 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D9_ACC_OUT</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>889.5,579,889.5,595.5</points>
<intersection>579 1</intersection>
<intersection>595.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>889.5,579,894.5,579</points>
<connection>
<GID>481</GID>
<name>IN_4</name></connection>
<intersection>889.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>889.5,595.5,891,595.5</points>
<connection>
<GID>742</GID>
<name>IN_0</name></connection>
<intersection>889.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>891,570.5,891,575</points>
<connection>
<GID>825</GID>
<name>IN_0</name></connection>
<intersection>575 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>891,575,894.5,575</points>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<intersection>891 0</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>890.5,567.5,890.5,576</points>
<intersection>567.5 2</intersection>
<intersection>576 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>890.5,576,894.5,576</points>
<connection>
<GID>481</GID>
<name>IN_1</name></connection>
<intersection>890.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>890.5,567.5,891,567.5</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<intersection>890.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>890,564.5,890,577</points>
<intersection>564.5 1</intersection>
<intersection>577 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>890,564.5,891,564.5</points>
<connection>
<GID>746</GID>
<name>IN_0</name></connection>
<intersection>890 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>890,577,894.5,577</points>
<connection>
<GID>481</GID>
<name>IN_2</name></connection>
<intersection>890 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>889.5,561.5,889.5,578</points>
<intersection>561.5 1</intersection>
<intersection>578 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>889.5,561.5,891,561.5</points>
<connection>
<GID>744</GID>
<name>IN_0</name></connection>
<intersection>889.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>889.5,578,894.5,578</points>
<connection>
<GID>481</GID>
<name>IN_3</name></connection>
<intersection>889.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>865.5,569.5,865.5,574.5</points>
<intersection>569.5 2</intersection>
<intersection>574.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>865.5,574.5,867,574.5</points>
<connection>
<GID>898</GID>
<name>IN_0</name></connection>
<intersection>865.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>865.5,569.5,867,569.5</points>
<connection>
<GID>841</GID>
<name>IN_0</name></connection>
<intersection>865.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>864.5,566.5,864.5,575.5</points>
<intersection>566.5 2</intersection>
<intersection>575.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>864.5,575.5,867,575.5</points>
<connection>
<GID>898</GID>
<name>IN_1</name></connection>
<intersection>864.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>864.5,566.5,867,566.5</points>
<connection>
<GID>842</GID>
<name>IN_0</name></connection>
<intersection>864.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>863.5,563.5,863.5,576.5</points>
<intersection>563.5 2</intersection>
<intersection>576.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>863.5,576.5,867,576.5</points>
<connection>
<GID>898</GID>
<name>IN_2</name></connection>
<intersection>863.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>863.5,563.5,867,563.5</points>
<connection>
<GID>843</GID>
<name>IN_0</name></connection>
<intersection>863.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>862.5,560.5,862.5,577.5</points>
<intersection>560.5 2</intersection>
<intersection>577.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>862.5,577.5,867,577.5</points>
<connection>
<GID>898</GID>
<name>IN_3</name></connection>
<intersection>862.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>862.5,560.5,867,560.5</points>
<connection>
<GID>844</GID>
<name>IN_0</name></connection>
<intersection>862.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>865.5,581.5,865.5,586.5</points>
<intersection>581.5 1</intersection>
<intersection>586.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>865.5,581.5,867,581.5</points>
<connection>
<GID>898</GID>
<name>IN_7</name></connection>
<intersection>865.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>865.5,586.5,867,586.5</points>
<connection>
<GID>850</GID>
<name>IN_0</name></connection>
<intersection>865.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>864.5,580.5,864.5,589.5</points>
<intersection>580.5 1</intersection>
<intersection>589.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>864.5,580.5,867,580.5</points>
<connection>
<GID>898</GID>
<name>IN_6</name></connection>
<intersection>864.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>864.5,589.5,867,589.5</points>
<connection>
<GID>848</GID>
<name>IN_0</name></connection>
<intersection>864.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>863.5,579.5,863.5,592.5</points>
<intersection>579.5 1</intersection>
<intersection>592.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>863.5,579.5,867,579.5</points>
<connection>
<GID>898</GID>
<name>IN_5</name></connection>
<intersection>863.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>863.5,592.5,867,592.5</points>
<connection>
<GID>846</GID>
<name>IN_0</name></connection>
<intersection>863.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>908,552.5,912,552.5</points>
<connection>
<GID>833</GID>
<name>OUT</name></connection>
<connection>
<GID>827</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>862.5,578.5,862.5,595.5</points>
<intersection>578.5 1</intersection>
<intersection>595.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>862.5,578.5,867,578.5</points>
<connection>
<GID>898</GID>
<name>IN_4</name></connection>
<intersection>862.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>862.5,595.5,867,595.5</points>
<connection>
<GID>845</GID>
<name>IN_0</name></connection>
<intersection>862.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>901.5,548.5,901.5,551.5</points>
<intersection>548.5 4</intersection>
<intersection>551.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>901.5,551.5,902,551.5</points>
<connection>
<GID>833</GID>
<name>IN_1</name></connection>
<intersection>901.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>901,548.5,901.5,548.5</points>
<connection>
<GID>832</GID>
<name>OUT</name></connection>
<intersection>901.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>892.5,546,892.5,547.5</points>
<intersection>546 2</intersection>
<intersection>547.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>892.5,547.5,895,547.5</points>
<connection>
<GID>832</GID>
<name>IN_1</name></connection>
<intersection>892.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>890.5,546,892.5,546</points>
<connection>
<GID>857</GID>
<name>CLK</name></connection>
<intersection>892.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>856,553.5,902,553.5</points>
<connection>
<GID>835</GID>
<name>OUT_0</name></connection>
<connection>
<GID>833</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>855.5,549,895,549</points>
<connection>
<GID>840</GID>
<name>OUT_0</name></connection>
<intersection>895 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>895,549,895,549.5</points>
<connection>
<GID>832</GID>
<name>IN_0</name></connection>
<intersection>549 1</intersection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>856,545.5,857.5,545.5</points>
<connection>
<GID>873</GID>
<name>IN_0</name></connection>
<connection>
<GID>870</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>912,582,912,586.5</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>582 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>912,582,915.5,582</points>
<connection>
<GID>281</GID>
<name>IN_7</name></connection>
<intersection>912 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>911.5,581,911.5,589.5</points>
<intersection>581 1</intersection>
<intersection>589.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>911.5,581,915.5,581</points>
<connection>
<GID>281</GID>
<name>IN_6</name></connection>
<intersection>911.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>911.5,589.5,912,589.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>911.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>911,580,911,592.5</points>
<intersection>580 1</intersection>
<intersection>592.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>911,580,915.5,580</points>
<connection>
<GID>281</GID>
<name>IN_5</name></connection>
<intersection>911 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>911,592.5,912,592.5</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>911 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>910.5,579,910.5,595.5</points>
<intersection>579 1</intersection>
<intersection>595.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>910.5,579,915.5,579</points>
<connection>
<GID>281</GID>
<name>IN_4</name></connection>
<intersection>910.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>910.5,595.5,912,595.5</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>910.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>912,570.5,912,575</points>
<connection>
<GID>460</GID>
<name>IN_0</name></connection>
<intersection>575 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>912,575,915.5,575</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>912 0</intersection></hsegment></shape></wire>
<wire>
<ID>679</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>850.5,569.5,850.5,574.5</points>
<intersection>569.5 1</intersection>
<intersection>574.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>850.5,569.5,851.5,569.5</points>
<connection>
<GID>859</GID>
<name>IN_0</name></connection>
<intersection>850.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>850.5,574.5,851.5,574.5</points>
<connection>
<GID>901</GID>
<name>IN_0</name></connection>
<intersection>850.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>680</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>849.5,566.5,849.5,575.5</points>
<intersection>566.5 2</intersection>
<intersection>575.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>849.5,575.5,851.5,575.5</points>
<connection>
<GID>901</GID>
<name>IN_1</name></connection>
<intersection>849.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>849.5,566.5,851.5,566.5</points>
<connection>
<GID>864</GID>
<name>IN_0</name></connection>
<intersection>849.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>681</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>848.5,563.5,848.5,576.5</points>
<intersection>563.5 2</intersection>
<intersection>576.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>848.5,576.5,851.5,576.5</points>
<connection>
<GID>901</GID>
<name>IN_2</name></connection>
<intersection>848.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>848.5,563.5,851.5,563.5</points>
<connection>
<GID>865</GID>
<name>IN_0</name></connection>
<intersection>848.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>682</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>847.5,560.5,847.5,577.5</points>
<intersection>560.5 2</intersection>
<intersection>577.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>847.5,577.5,851.5,577.5</points>
<connection>
<GID>901</GID>
<name>IN_3</name></connection>
<intersection>847.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>847.5,560.5,851.5,560.5</points>
<connection>
<GID>867</GID>
<name>IN_0</name></connection>
<intersection>847.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>683</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>827.5,570.5,827.5,575</points>
<intersection>570.5 2</intersection>
<intersection>575 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>827.5,575,828.5,575</points>
<connection>
<GID>893</GID>
<name>IN_0</name></connection>
<intersection>827.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>827.5,570.5,828.5,570.5</points>
<connection>
<GID>899</GID>
<name>IN_0</name></connection>
<intersection>827.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>684</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>826.5,567.5,826.5,576</points>
<intersection>567.5 2</intersection>
<intersection>576 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>826.5,576,828.5,576</points>
<connection>
<GID>893</GID>
<name>IN_1</name></connection>
<intersection>826.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>826.5,567.5,828.5,567.5</points>
<connection>
<GID>900</GID>
<name>IN_0</name></connection>
<intersection>826.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>685</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>825.5,564.5,825.5,577</points>
<intersection>564.5 2</intersection>
<intersection>577 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>825.5,577,828.5,577</points>
<connection>
<GID>893</GID>
<name>IN_2</name></connection>
<intersection>825.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>825.5,564.5,828.5,564.5</points>
<connection>
<GID>902</GID>
<name>IN_0</name></connection>
<intersection>825.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>689</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>824.5,561.5,824.5,578</points>
<intersection>561.5 2</intersection>
<intersection>578 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>824.5,578,828.5,578</points>
<connection>
<GID>893</GID>
<name>IN_3</name></connection>
<intersection>824.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>824.5,561.5,828.5,561.5</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>824.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>911.5,567.5,911.5,576</points>
<intersection>567.5 2</intersection>
<intersection>576 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>911.5,576,915.5,576</points>
<connection>
<GID>281</GID>
<name>IN_1</name></connection>
<intersection>911.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>911.5,567.5,912,567.5</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<intersection>911.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>911,564.5,911,577</points>
<intersection>564.5 1</intersection>
<intersection>577 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>911,564.5,912,564.5</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>911 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>911,577,915.5,577</points>
<connection>
<GID>281</GID>
<name>IN_2</name></connection>
<intersection>911 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>910.5,561.5,910.5,578</points>
<intersection>561.5 1</intersection>
<intersection>578 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>910.5,561.5,912,561.5</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>910.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>910.5,578,915.5,578</points>
<connection>
<GID>281</GID>
<name>IN_3</name></connection>
<intersection>910.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>891,582,891,586.5</points>
<connection>
<GID>736</GID>
<name>IN_0</name></connection>
<intersection>582 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>891,582,894.5,582</points>
<connection>
<GID>481</GID>
<name>IN_7</name></connection>
<intersection>891 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>890.5,581,890.5,589.5</points>
<intersection>581 1</intersection>
<intersection>589.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>890.5,581,894.5,581</points>
<connection>
<GID>481</GID>
<name>IN_6</name></connection>
<intersection>890.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>890.5,589.5,891,589.5</points>
<connection>
<GID>738</GID>
<name>IN_0</name></connection>
<intersection>890.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>890,580,890,592.5</points>
<intersection>580 1</intersection>
<intersection>592.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>890,580,894.5,580</points>
<connection>
<GID>481</GID>
<name>IN_5</name></connection>
<intersection>890 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>890,592.5,891,592.5</points>
<connection>
<GID>740</GID>
<name>IN_0</name></connection>
<intersection>890 0</intersection></hsegment></shape></wire></page 8>
<page 9>
<PageViewport>757.886,1092.07,966.952,984.247</PageViewport>
<gate>
<ID>272</ID>
<type>DA_FROM</type>
<position>807.5,1041.5</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA3</lparam></gate>
<gate>
<ID>278</ID>
<type>DA_FROM</type>
<position>807.5,1044.5</position>
<input>
<ID>IN_0</ID>690 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA4</lparam></gate>
<gate>
<ID>290</ID>
<type>DA_FROM</type>
<position>807.5,1047.5</position>
<input>
<ID>IN_0</ID>691 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA5</lparam></gate>
<gate>
<ID>297</ID>
<type>DA_FROM</type>
<position>807.5,1050.5</position>
<input>
<ID>IN_0</ID>692 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA6</lparam></gate>
<gate>
<ID>106</ID>
<type>DE_TO</type>
<position>862,1027.5</position>
<input>
<ID>IN_0</ID>716 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD5</lparam></gate>
<gate>
<ID>110</ID>
<type>DE_TO</type>
<position>862,1024.5</position>
<input>
<ID>IN_0</ID>717 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD6</lparam></gate>
<gate>
<ID>111</ID>
<type>DE_TO</type>
<position>862,1021.5</position>
<input>
<ID>IN_0</ID>718 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD7</lparam></gate>
<gate>
<ID>112</ID>
<type>DE_TO</type>
<position>862,1003.5</position>
<input>
<ID>IN_0</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD13</lparam></gate>
<gate>
<ID>114</ID>
<type>DE_TO</type>
<position>862,1000.5</position>
<input>
<ID>IN_0</ID>731 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD14</lparam></gate>
<gate>
<ID>308</ID>
<type>DA_FROM</type>
<position>807.5,1053.5</position>
<input>
<ID>IN_0</ID>693 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA7</lparam></gate>
<gate>
<ID>115</ID>
<type>DE_TO</type>
<position>862,997.5</position>
<input>
<ID>IN_0</ID>732 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD15</lparam></gate>
<gate>
<ID>116</ID>
<type>DE_TO</type>
<position>862,1018.5</position>
<input>
<ID>IN_0</ID>719 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD8</lparam></gate>
<gate>
<ID>117</ID>
<type>DE_TO</type>
<position>862,1015.5</position>
<input>
<ID>IN_0</ID>720 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD9</lparam></gate>
<gate>
<ID>118</ID>
<type>DE_TO</type>
<position>862,1012.5</position>
<input>
<ID>IN_0</ID>724 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD10</lparam></gate>
<gate>
<ID>119</ID>
<type>DE_TO</type>
<position>862,1009.5</position>
<input>
<ID>IN_0</ID>728 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD11</lparam></gate>
<gate>
<ID>120</ID>
<type>DE_TO</type>
<position>862,1006.5</position>
<input>
<ID>IN_0</ID>729 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD12</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>831,1078</position>
<gparam>LABEL_TEXT Memoria de Programa</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>BI_ROM_12x16</type>
<position>843.5,1054</position>
<input>
<ID>ADDRESS_0</ID>57 </input>
<input>
<ID>ADDRESS_1</ID>58 </input>
<input>
<ID>ADDRESS_10</ID>708 </input>
<input>
<ID>ADDRESS_11</ID>709 </input>
<input>
<ID>ADDRESS_2</ID>59 </input>
<input>
<ID>ADDRESS_3</ID>72 </input>
<input>
<ID>ADDRESS_4</ID>690 </input>
<input>
<ID>ADDRESS_5</ID>691 </input>
<input>
<ID>ADDRESS_6</ID>692 </input>
<input>
<ID>ADDRESS_7</ID>693 </input>
<input>
<ID>ADDRESS_8</ID>700 </input>
<input>
<ID>ADDRESS_9</ID>701 </input>
<output>
<ID>DATA_OUT_0</ID>711 </output>
<output>
<ID>DATA_OUT_1</ID>712 </output>
<output>
<ID>DATA_OUT_10</ID>724 </output>
<output>
<ID>DATA_OUT_11</ID>728 </output>
<output>
<ID>DATA_OUT_12</ID>729 </output>
<output>
<ID>DATA_OUT_13</ID>730 </output>
<output>
<ID>DATA_OUT_14</ID>731 </output>
<output>
<ID>DATA_OUT_15</ID>732 </output>
<output>
<ID>DATA_OUT_2</ID>713 </output>
<output>
<ID>DATA_OUT_3</ID>714 </output>
<output>
<ID>DATA_OUT_4</ID>715 </output>
<output>
<ID>DATA_OUT_5</ID>716 </output>
<output>
<ID>DATA_OUT_6</ID>717 </output>
<output>
<ID>DATA_OUT_7</ID>718 </output>
<output>
<ID>DATA_OUT_8</ID>719 </output>
<output>
<ID>DATA_OUT_9</ID>720 </output>
<input>
<ID>ENABLE_0</ID>710 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:0 32770</lparam>
<lparam>Address:1 32776</lparam>
<lparam>Address:2 8191</lparam>
<lparam>Address:3 10922</lparam>
<lparam>Address:4 13395</lparam>
<lparam>Address:5 36864</lparam>
<lparam>Address:6 32769</lparam>
<lparam>Address:8 17491</lparam>
<lparam>Address:9 21587</lparam>
<lparam>Address:10 25683</lparam>
<lparam>Address:11 29779</lparam>
<lparam>Address:12 5203</lparam>
<lparam>Address:13 9299</lparam>
<lparam>Address:14 13395</lparam>
<lparam>Address:15 17491</lparam>
<lparam>Address:16 21587</lparam>
<lparam>Address:17 25683</lparam>
<lparam>Address:18 29779</lparam>
<lparam>Address:19 5203</lparam>
<lparam>Address:20 9299</lparam>
<lparam>Address:21 13395</lparam>
<lparam>Address:22 17491</lparam>
<lparam>Address:23 21587</lparam>
<lparam>Address:24 25683</lparam>
<lparam>Address:25 29779</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>807.5,1032.5</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA0</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>807.5,1035.5</position>
<input>
<ID>IN_0</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA1</lparam></gate>
<gate>
<ID>906</ID>
<type>DA_FROM</type>
<position>807.5,1056.5</position>
<input>
<ID>IN_0</ID>700 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA8</lparam></gate>
<gate>
<ID>134</ID>
<type>DA_FROM</type>
<position>807.5,1038.5</position>
<input>
<ID>IN_0</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA2</lparam></gate>
<gate>
<ID>907</ID>
<type>DA_FROM</type>
<position>807.5,1059.5</position>
<input>
<ID>IN_0</ID>701 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA9</lparam></gate>
<gate>
<ID>908</ID>
<type>DA_FROM</type>
<position>807.5,1062.5</position>
<input>
<ID>IN_0</ID>708 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA10</lparam></gate>
<gate>
<ID>909</ID>
<type>DA_FROM</type>
<position>807.5,1065.5</position>
<input>
<ID>IN_0</ID>709 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCA11</lparam></gate>
<gate>
<ID>910</ID>
<type>EE_VDD</type>
<position>854,1055.5</position>
<output>
<ID>OUT_0</ID>710 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>911</ID>
<type>DE_TO</type>
<position>862,1042.5</position>
<input>
<ID>IN_0</ID>711 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD0</lparam></gate>
<gate>
<ID>912</ID>
<type>DE_TO</type>
<position>862,1039.5</position>
<input>
<ID>IN_0</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD1</lparam></gate>
<gate>
<ID>913</ID>
<type>DE_TO</type>
<position>862,1036.5</position>
<input>
<ID>IN_0</ID>713 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD2</lparam></gate>
<gate>
<ID>914</ID>
<type>DE_TO</type>
<position>862,1033.5</position>
<input>
<ID>IN_0</ID>714 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD3</lparam></gate>
<gate>
<ID>915</ID>
<type>DE_TO</type>
<position>862,1030.5</position>
<input>
<ID>IN_0</ID>715 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PD4</lparam></gate>
<gate>
<ID>916</ID>
<type>AA_LABEL</type>
<position>830.5,1087.5</position>
<gparam>LABEL_TEXT Prof.  Angelo Zanini / Nuncio Perrella</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>923</ID>
<type>AA_LABEL</type>
<position>836,1099</position>
<gparam>LABEL_TEXT PROCESSADOR BIP IMT - MAUA 2022</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0</gparam></gate>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>833,1032.5,833,1048.5</points>
<intersection>1032.5 2</intersection>
<intersection>1048.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>833,1048.5,834.5,1048.5</points>
<connection>
<GID>122</GID>
<name>ADDRESS_0</name></connection>
<intersection>833 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>809.5,1032.5,833,1032.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>833 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>832,1035.5,832,1049.5</points>
<intersection>1035.5 2</intersection>
<intersection>1049.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>832,1049.5,834.5,1049.5</points>
<connection>
<GID>122</GID>
<name>ADDRESS_1</name></connection>
<intersection>832 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>809.5,1035.5,832,1035.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>832 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>831,1038.5,831,1050.5</points>
<intersection>1038.5 2</intersection>
<intersection>1050.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>831,1050.5,834.5,1050.5</points>
<connection>
<GID>122</GID>
<name>ADDRESS_2</name></connection>
<intersection>831 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>809.5,1038.5,831,1038.5</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>831 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>830,1041.5,830,1051.5</points>
<intersection>1041.5 2</intersection>
<intersection>1051.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>830,1051.5,834.5,1051.5</points>
<connection>
<GID>122</GID>
<name>ADDRESS_3</name></connection>
<intersection>830 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>809.5,1041.5,830,1041.5</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>830 0</intersection></hsegment></shape></wire>
<wire>
<ID>690</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>829,1044.5,829,1052.5</points>
<intersection>1044.5 2</intersection>
<intersection>1052.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>829,1052.5,834.5,1052.5</points>
<connection>
<GID>122</GID>
<name>ADDRESS_4</name></connection>
<intersection>829 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>809.5,1044.5,829,1044.5</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>829 0</intersection></hsegment></shape></wire>
<wire>
<ID>691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>828,1047.5,828,1053.5</points>
<intersection>1047.5 2</intersection>
<intersection>1053.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>828,1053.5,834.5,1053.5</points>
<connection>
<GID>122</GID>
<name>ADDRESS_5</name></connection>
<intersection>828 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>809.5,1047.5,828,1047.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>828 0</intersection></hsegment></shape></wire>
<wire>
<ID>692</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>827,1050.5,827,1054.5</points>
<intersection>1050.5 2</intersection>
<intersection>1054.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>827,1054.5,834.5,1054.5</points>
<connection>
<GID>122</GID>
<name>ADDRESS_6</name></connection>
<intersection>827 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>809.5,1050.5,827,1050.5</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>827 0</intersection></hsegment></shape></wire>
<wire>
<ID>693</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>826,1053.5,826,1055.5</points>
<intersection>1053.5 2</intersection>
<intersection>1055.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>826,1055.5,834.5,1055.5</points>
<connection>
<GID>122</GID>
<name>ADDRESS_7</name></connection>
<intersection>826 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>809.5,1053.5,826,1053.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>826 0</intersection></hsegment></shape></wire>
<wire>
<ID>700</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>809.5,1056.5,834.5,1056.5</points>
<connection>
<GID>906</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>ADDRESS_8</name></connection></hsegment></shape></wire>
<wire>
<ID>701</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>826,1057.5,826,1059.5</points>
<intersection>1057.5 1</intersection>
<intersection>1059.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>826,1057.5,834.5,1057.5</points>
<connection>
<GID>122</GID>
<name>ADDRESS_9</name></connection>
<intersection>826 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>809.5,1059.5,826,1059.5</points>
<connection>
<GID>907</GID>
<name>IN_0</name></connection>
<intersection>826 0</intersection></hsegment></shape></wire>
<wire>
<ID>708</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>827,1058.5,827,1062.5</points>
<intersection>1058.5 1</intersection>
<intersection>1062.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>827,1058.5,834.5,1058.5</points>
<connection>
<GID>122</GID>
<name>ADDRESS_10</name></connection>
<intersection>827 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>809.5,1062.5,827,1062.5</points>
<connection>
<GID>908</GID>
<name>IN_0</name></connection>
<intersection>827 0</intersection></hsegment></shape></wire>
<wire>
<ID>709</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>828,1059.5,828,1065.5</points>
<intersection>1059.5 1</intersection>
<intersection>1065.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>828,1059.5,834.5,1059.5</points>
<connection>
<GID>122</GID>
<name>ADDRESS_11</name></connection>
<intersection>828 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>809.5,1065.5,828,1065.5</points>
<connection>
<GID>909</GID>
<name>IN_0</name></connection>
<intersection>828 0</intersection></hsegment></shape></wire>
<wire>
<ID>710</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>852.5,1053.5,854,1053.5</points>
<connection>
<GID>122</GID>
<name>ENABLE_0</name></connection>
<intersection>854 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>854,1053.5,854,1054.5</points>
<connection>
<GID>910</GID>
<name>OUT_0</name></connection>
<intersection>1053.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>711</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>851,1042.5,860,1042.5</points>
<connection>
<GID>911</GID>
<name>IN_0</name></connection>
<intersection>851 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>851,1042.5,851,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_0</name></connection>
<intersection>1042.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>712</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>850,1039.5,850,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_1</name></connection>
<intersection>1039.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>850,1039.5,860,1039.5</points>
<connection>
<GID>912</GID>
<name>IN_0</name></connection>
<intersection>850 0</intersection></hsegment></shape></wire>
<wire>
<ID>713</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>849,1036.5,849,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_2</name></connection>
<intersection>1036.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>849,1036.5,860,1036.5</points>
<connection>
<GID>913</GID>
<name>IN_0</name></connection>
<intersection>849 0</intersection></hsegment></shape></wire>
<wire>
<ID>714</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>848,1033.5,848,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_3</name></connection>
<intersection>1033.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>848,1033.5,860,1033.5</points>
<connection>
<GID>914</GID>
<name>IN_0</name></connection>
<intersection>848 0</intersection></hsegment></shape></wire>
<wire>
<ID>715</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>847,1030.5,847,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_4</name></connection>
<intersection>1030.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>847,1030.5,860,1030.5</points>
<connection>
<GID>915</GID>
<name>IN_0</name></connection>
<intersection>847 0</intersection></hsegment></shape></wire>
<wire>
<ID>716</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>846,1027.5,846,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_5</name></connection>
<intersection>1027.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>846,1027.5,860,1027.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>846 0</intersection></hsegment></shape></wire>
<wire>
<ID>717</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>845,1024.5,845,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_6</name></connection>
<intersection>1024.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>845,1024.5,860,1024.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>845 0</intersection></hsegment></shape></wire>
<wire>
<ID>718</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>844,1021.5,844,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_7</name></connection>
<intersection>1021.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>844,1021.5,860,1021.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>844 0</intersection></hsegment></shape></wire>
<wire>
<ID>719</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>843,1018.5,843,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_8</name></connection>
<intersection>1018.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>843,1018.5,860,1018.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>843 0</intersection></hsegment></shape></wire>
<wire>
<ID>720</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>842,1015.5,842,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_9</name></connection>
<intersection>1015.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>842,1015.5,860,1015.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>842 0</intersection></hsegment></shape></wire>
<wire>
<ID>724</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>841,1012.5,841,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_10</name></connection>
<intersection>1012.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>841,1012.5,860,1012.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>841 0</intersection></hsegment></shape></wire>
<wire>
<ID>728</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>840,1009.5,840,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_11</name></connection>
<intersection>1009.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>840,1009.5,860,1009.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>840 0</intersection></hsegment></shape></wire>
<wire>
<ID>729</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>839,1006.5,839,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_12</name></connection>
<intersection>1006.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>839,1006.5,860,1006.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>839 0</intersection></hsegment></shape></wire>
<wire>
<ID>730</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>838,1003.5,838,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_13</name></connection>
<intersection>1003.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>838,1003.5,860,1003.5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>838 0</intersection></hsegment></shape></wire>
<wire>
<ID>731</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>837,1000.5,837,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_14</name></connection>
<intersection>1000.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>837,1000.5,860,1000.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>837 0</intersection></hsegment></shape></wire>
<wire>
<ID>732</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>836,997.5,836,1043</points>
<connection>
<GID>122</GID>
<name>DATA_OUT_15</name></connection>
<intersection>997.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>836,997.5,860,997.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>836 0</intersection></hsegment></shape></wire></page 9></circuit>